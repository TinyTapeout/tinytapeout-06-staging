VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_openframe_mask_rev
  CLASS BLOCK ;
  FOREIGN tt_um_openframe_mask_rev ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.910 2.480 41.510 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.860 2.480 79.460 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.810 2.480 117.410 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.760 2.480 155.360 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.935 2.480 22.535 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.885 2.480 60.485 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.835 2.480 98.435 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.785 2.480 136.385 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 110.520 134.930 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END ena
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 21.470 0.000 21.770 1.000 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 49.070 0.000 49.370 1.000 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 0.000 52.130 1.000 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 54.590 0.000 54.890 1.000 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 57.350 0.000 57.650 1.000 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 60.110 0.000 60.410 1.000 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 0.000 63.170 1.000 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 65.630 0.000 65.930 1.000 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 68.390 0.000 68.690 1.000 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 71.150 0.000 71.450 1.000 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 73.910 0.000 74.210 1.000 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 24.230 0.000 24.530 1.000 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 76.670 0.000 76.970 1.000 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 79.430 0.000 79.730 1.000 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 82.190 0.000 82.490 1.000 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 0.000 85.250 1.000 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 87.710 0.000 88.010 1.000 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 90.470 0.000 90.770 1.000 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 93.230 0.000 93.530 1.000 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 95.990 0.000 96.290 1.000 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 98.750 0.000 99.050 1.000 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 101.510 0.000 101.810 1.000 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 26.990 0.000 27.290 1.000 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 104.270 0.000 104.570 1.000 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 0.000 107.330 1.000 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 0.000 30.050 1.000 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 32.510 0.000 32.810 1.000 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 35.270 0.000 35.570 1.000 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 38.030 0.000 38.330 1.000 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 0.000 41.090 1.000 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 43.550 0.000 43.850 1.000 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 46.310 0.000 46.610 1.000 ;
    END
  END mask_rev[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 123.590 110.520 123.890 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.550 110.520 112.850 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 110.520 101.810 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.470 110.520 90.770 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.710 110.520 88.010 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.270 110.520 35.570 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 110.520 30.050 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.230 110.520 24.530 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 62.870 110.520 63.170 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 60.110 110.520 60.410 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 57.350 110.520 57.650 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 54.590 110.520 54.890 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.520 52.130 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 49.070 110.520 49.370 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 46.310 110.520 46.610 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 43.550 110.520 43.850 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 110.520 85.250 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER met4 ;
        RECT 82.190 110.520 82.490 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 79.430 110.520 79.730 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 76.670 110.520 76.970 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.933750 ;
    PORT
      LAYER met4 ;
        RECT 73.910 110.520 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 71.150 110.520 71.450 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 68.390 110.520 68.690 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.630 110.520 65.930 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 154.750 108.990 ;
        RECT 2.570 101.945 154.750 104.775 ;
        RECT 2.570 96.505 154.750 99.335 ;
        RECT 2.570 91.065 154.750 93.895 ;
        RECT 2.570 85.625 154.750 88.455 ;
        RECT 2.570 80.185 154.750 83.015 ;
        RECT 2.570 74.745 154.750 77.575 ;
        RECT 2.570 69.305 154.750 72.135 ;
        RECT 2.570 63.865 154.750 66.695 ;
        RECT 2.570 58.425 154.750 61.255 ;
        RECT 2.570 52.985 154.750 55.815 ;
        RECT 2.570 47.545 154.750 50.375 ;
        RECT 2.570 42.105 154.750 44.935 ;
        RECT 2.570 36.665 154.750 39.495 ;
        RECT 2.570 31.225 154.750 34.055 ;
        RECT 2.570 25.785 154.750 28.615 ;
        RECT 2.570 20.345 154.750 23.175 ;
        RECT 2.570 14.905 154.750 17.735 ;
        RECT 2.570 9.465 154.750 12.295 ;
        RECT 2.570 4.025 154.750 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 154.560 108.885 ;
      LAYER met1 ;
        RECT 2.760 0.040 155.360 109.040 ;
      LAYER met2 ;
        RECT 20.965 0.010 155.330 110.005 ;
      LAYER met3 ;
        RECT 20.945 0.175 155.350 109.985 ;
      LAYER met4 ;
        RECT 22.170 110.120 23.830 111.170 ;
        RECT 24.930 110.120 26.590 111.170 ;
        RECT 27.690 110.120 29.350 111.170 ;
        RECT 30.450 110.120 32.110 111.170 ;
        RECT 33.210 110.120 34.870 111.170 ;
        RECT 35.970 110.120 37.630 111.170 ;
        RECT 38.730 110.120 40.390 111.170 ;
        RECT 41.490 110.120 43.150 111.170 ;
        RECT 44.250 110.120 45.910 111.170 ;
        RECT 47.010 110.120 48.670 111.170 ;
        RECT 49.770 110.120 51.430 111.170 ;
        RECT 52.530 110.120 54.190 111.170 ;
        RECT 55.290 110.120 56.950 111.170 ;
        RECT 58.050 110.120 59.710 111.170 ;
        RECT 60.810 110.120 62.470 111.170 ;
        RECT 63.570 110.120 65.230 111.170 ;
        RECT 66.330 110.120 67.990 111.170 ;
        RECT 69.090 110.120 70.750 111.170 ;
        RECT 71.850 110.120 73.510 111.170 ;
        RECT 74.610 110.120 76.270 111.170 ;
        RECT 77.370 110.120 79.030 111.170 ;
        RECT 80.130 110.120 81.790 111.170 ;
        RECT 82.890 110.120 84.550 111.170 ;
        RECT 85.650 110.120 87.310 111.170 ;
        RECT 88.410 110.120 90.070 111.170 ;
        RECT 91.170 110.120 92.830 111.170 ;
        RECT 93.930 110.120 95.590 111.170 ;
        RECT 96.690 110.120 98.350 111.170 ;
        RECT 99.450 110.120 101.110 111.170 ;
        RECT 102.210 110.120 103.870 111.170 ;
        RECT 104.970 110.120 106.630 111.170 ;
        RECT 107.730 110.120 109.390 111.170 ;
        RECT 110.490 110.120 112.150 111.170 ;
        RECT 113.250 110.120 114.910 111.170 ;
        RECT 116.010 110.120 117.670 111.170 ;
        RECT 118.770 110.120 120.430 111.170 ;
        RECT 121.530 110.120 123.190 111.170 ;
        RECT 124.290 110.120 125.950 111.170 ;
        RECT 127.050 110.120 128.710 111.170 ;
        RECT 21.455 109.440 129.425 110.120 ;
        RECT 22.935 2.080 39.510 109.440 ;
        RECT 41.910 2.080 58.485 109.440 ;
        RECT 60.885 2.080 77.460 109.440 ;
        RECT 79.860 2.080 96.435 109.440 ;
        RECT 98.835 2.080 115.410 109.440 ;
        RECT 117.810 2.080 129.425 109.440 ;
        RECT 21.455 1.400 129.425 2.080 ;
        RECT 22.170 0.175 23.830 1.400 ;
        RECT 24.930 0.175 26.590 1.400 ;
        RECT 27.690 0.175 29.350 1.400 ;
        RECT 30.450 0.175 32.110 1.400 ;
        RECT 33.210 0.175 34.870 1.400 ;
        RECT 35.970 0.175 37.630 1.400 ;
        RECT 38.730 0.175 40.390 1.400 ;
        RECT 41.490 0.175 43.150 1.400 ;
        RECT 44.250 0.175 45.910 1.400 ;
        RECT 47.010 0.175 48.670 1.400 ;
        RECT 49.770 0.175 51.430 1.400 ;
        RECT 52.530 0.175 54.190 1.400 ;
        RECT 55.290 0.175 56.950 1.400 ;
        RECT 58.050 0.175 59.710 1.400 ;
        RECT 60.810 0.175 62.470 1.400 ;
        RECT 63.570 0.175 65.230 1.400 ;
        RECT 66.330 0.175 67.990 1.400 ;
        RECT 69.090 0.175 70.750 1.400 ;
        RECT 71.850 0.175 73.510 1.400 ;
        RECT 74.610 0.175 76.270 1.400 ;
        RECT 77.370 0.175 79.030 1.400 ;
        RECT 80.130 0.175 81.790 1.400 ;
        RECT 82.890 0.175 84.550 1.400 ;
        RECT 85.650 0.175 87.310 1.400 ;
        RECT 88.410 0.175 90.070 1.400 ;
        RECT 91.170 0.175 92.830 1.400 ;
        RECT 93.930 0.175 95.590 1.400 ;
        RECT 96.690 0.175 98.350 1.400 ;
        RECT 99.450 0.175 101.110 1.400 ;
        RECT 102.210 0.175 103.870 1.400 ;
        RECT 104.970 0.175 106.630 1.400 ;
        RECT 107.730 0.175 129.425 1.400 ;
  END
END tt_um_openframe_mask_rev
END LIBRARY

