VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_r2r_dac
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_r2r_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 0.000 2.500 225.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 0.000 50.500 225.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 110.980 106.360 111.310 106.530 ;
        RECT 112.590 106.400 112.920 106.570 ;
        RECT 111.060 104.545 111.230 106.360 ;
        RECT 112.670 104.585 112.840 106.400 ;
        RECT 114.410 106.380 114.740 106.550 ;
        RECT 114.490 104.565 114.660 106.380 ;
        RECT 116.080 106.320 116.410 106.490 ;
        RECT 118.100 106.340 118.430 106.510 ;
        RECT 116.160 104.505 116.330 106.320 ;
        RECT 118.180 104.525 118.350 106.340 ;
        RECT 111.060 88.870 111.230 90.685 ;
        RECT 112.670 88.910 112.840 90.725 ;
        RECT 110.980 88.700 111.310 88.870 ;
        RECT 112.590 88.740 112.920 88.910 ;
        RECT 114.490 88.890 114.660 90.705 ;
        RECT 114.410 88.720 114.740 88.890 ;
        RECT 116.160 88.830 116.330 90.645 ;
        RECT 118.180 88.850 118.350 90.665 ;
        RECT 116.080 88.660 116.410 88.830 ;
        RECT 118.100 88.680 118.430 88.850 ;
        RECT 112.840 87.150 113.170 87.320 ;
        RECT 112.920 85.335 113.090 87.150 ;
        RECT 115.040 87.140 115.370 87.310 ;
        RECT 117.200 87.210 117.530 87.380 ;
        RECT 115.120 85.325 115.290 87.140 ;
        RECT 117.280 85.395 117.450 87.210 ;
        RECT 112.920 76.500 113.090 78.315 ;
        RECT 112.840 76.330 113.170 76.500 ;
        RECT 115.120 76.490 115.290 78.305 ;
        RECT 117.280 76.560 117.450 78.375 ;
        RECT 115.040 76.320 115.370 76.490 ;
        RECT 117.200 76.390 117.530 76.560 ;
      LAYER mcon ;
        RECT 111.060 88.700 111.230 90.685 ;
        RECT 112.670 88.740 112.840 90.725 ;
        RECT 114.490 88.720 114.660 90.705 ;
        RECT 116.160 88.660 116.330 90.645 ;
        RECT 118.180 88.680 118.350 90.665 ;
        RECT 112.920 76.330 113.090 78.315 ;
        RECT 115.120 76.320 115.290 78.305 ;
        RECT 117.280 76.390 117.450 78.375 ;
      LAYER met1 ;
        RECT 110.540 112.470 111.310 113.030 ;
        RECT 112.490 112.500 113.260 113.060 ;
        RECT 115.660 112.560 116.430 113.120 ;
        RECT 118.850 112.560 119.620 113.120 ;
        RECT 110.600 110.040 111.020 112.470 ;
        RECT 112.640 110.660 113.060 112.500 ;
        RECT 115.790 111.130 116.210 112.560 ;
        RECT 115.790 110.710 116.490 111.130 ;
        RECT 112.640 110.240 114.860 110.660 ;
        RECT 110.600 109.620 112.980 110.040 ;
        RECT 111.030 106.555 111.260 106.590 ;
        RECT 106.960 105.965 111.435 106.555 ;
        RECT 112.560 105.990 112.980 109.620 ;
        RECT 114.440 105.990 114.860 110.240 ;
        RECT 105.240 105.100 106.570 105.450 ;
        RECT 106.960 105.100 107.550 105.965 ;
        RECT 105.240 104.510 107.550 105.100 ;
        RECT 105.240 104.240 106.570 104.510 ;
        RECT 111.030 104.485 111.260 105.965 ;
        RECT 112.640 104.525 112.870 105.990 ;
        RECT 114.460 104.505 114.690 105.990 ;
        RECT 116.070 105.980 116.490 110.710 ;
        RECT 119.020 108.820 119.440 112.560 ;
        RECT 118.090 108.400 119.440 108.820 ;
        RECT 118.090 106.020 118.510 108.400 ;
        RECT 116.130 104.445 116.360 105.980 ;
        RECT 118.150 104.465 118.380 106.020 ;
        RECT 111.030 90.590 111.260 90.745 ;
        RECT 112.640 90.590 112.870 90.785 ;
        RECT 110.700 88.670 113.070 90.590 ;
        RECT 114.460 89.350 114.690 90.765 ;
        RECT 114.370 89.255 114.800 89.350 ;
        RECT 116.130 89.310 116.360 90.705 ;
        RECT 118.150 89.310 118.380 90.725 ;
        RECT 116.030 89.265 116.460 89.310 ;
        RECT 111.030 88.640 111.665 88.670 ;
        RECT 111.140 75.945 111.665 88.640 ;
        RECT 114.370 88.610 114.805 89.255 ;
        RECT 114.375 88.265 114.805 88.610 ;
        RECT 112.790 87.835 114.805 88.265 ;
        RECT 116.025 88.570 116.460 89.265 ;
        RECT 118.070 89.295 118.500 89.310 ;
        RECT 118.070 88.570 118.525 89.295 ;
        RECT 128.920 88.940 129.580 89.440 ;
        RECT 112.790 86.920 113.220 87.835 ;
        RECT 112.890 85.275 113.120 86.920 ;
        RECT 112.890 77.070 113.120 78.375 ;
        RECT 112.760 75.945 113.250 77.070 ;
        RECT 113.645 76.695 114.075 87.835 ;
        RECT 116.025 87.770 116.455 88.570 ;
        RECT 118.095 87.825 118.525 88.570 ;
        RECT 128.935 87.825 129.365 88.940 ;
        RECT 118.095 87.780 129.365 87.825 ;
        RECT 115.020 87.340 116.455 87.770 ;
        RECT 115.020 87.030 115.450 87.340 ;
        RECT 115.090 85.265 115.320 87.030 ;
        RECT 115.090 76.695 115.320 78.365 ;
        RECT 113.645 76.265 115.505 76.695 ;
        RECT 116.025 76.655 116.455 87.340 ;
        RECT 117.190 87.395 129.365 87.780 ;
        RECT 117.190 87.350 118.525 87.395 ;
        RECT 117.190 87.040 117.620 87.350 ;
        RECT 117.250 85.335 117.480 87.040 ;
        RECT 117.250 76.655 117.480 78.435 ;
        RECT 115.090 76.260 115.320 76.265 ;
        RECT 116.025 76.225 117.535 76.655 ;
        RECT 111.140 75.455 113.250 75.945 ;
        RECT 111.140 75.440 111.665 75.455 ;
      LAYER via ;
        RECT 110.590 112.470 111.260 113.030 ;
        RECT 112.540 112.500 113.210 113.060 ;
        RECT 115.710 112.560 116.380 113.120 ;
        RECT 118.900 112.560 119.570 113.120 ;
        RECT 105.290 104.240 106.520 105.450 ;
        RECT 128.970 88.940 129.530 89.440 ;
      LAYER met2 ;
        RECT 110.590 112.420 111.260 113.080 ;
        RECT 112.540 112.450 113.210 113.110 ;
        RECT 115.710 112.510 116.380 113.170 ;
        RECT 118.900 112.510 119.570 113.170 ;
        RECT 105.290 104.190 106.520 105.500 ;
        RECT 128.970 88.890 129.530 89.490 ;
      LAYER via2 ;
        RECT 110.590 112.470 111.260 113.030 ;
        RECT 112.540 112.500 113.210 113.060 ;
        RECT 115.710 112.560 116.380 113.120 ;
        RECT 118.900 112.560 119.570 113.120 ;
        RECT 105.290 104.240 106.520 105.450 ;
        RECT 128.970 88.940 129.530 89.440 ;
      LAYER met3 ;
        RECT 110.540 112.445 111.310 113.055 ;
        RECT 112.490 112.475 113.260 113.085 ;
        RECT 115.660 112.535 116.430 113.145 ;
        RECT 118.850 112.535 119.620 113.145 ;
        RECT 105.240 104.215 106.570 105.475 ;
        RECT 128.920 88.915 129.580 89.465 ;
      LAYER via3 ;
        RECT 110.590 112.470 111.260 113.030 ;
        RECT 112.540 112.500 113.210 113.060 ;
        RECT 115.710 112.560 116.380 113.120 ;
        RECT 118.900 112.560 119.570 113.120 ;
        RECT 105.290 104.240 106.520 105.450 ;
        RECT 128.970 88.940 129.530 89.440 ;
      LAYER met4 ;
        RECT 136.470 133.810 136.770 224.760 ;
        RECT 110.750 133.510 136.770 133.810 ;
        RECT 110.750 113.035 111.050 133.510 ;
        RECT 140.150 130.460 140.450 224.760 ;
        RECT 112.750 130.160 140.450 130.460 ;
        RECT 112.750 113.065 113.050 130.160 ;
        RECT 143.830 126.870 144.130 224.760 ;
        RECT 115.910 126.570 144.130 126.870 ;
        RECT 115.910 113.125 116.210 126.570 ;
        RECT 147.510 124.410 147.810 224.760 ;
        RECT 119.070 124.110 147.810 124.410 ;
        RECT 119.070 113.125 119.370 124.110 ;
        RECT 110.585 112.465 111.265 113.035 ;
        RECT 112.535 112.495 113.215 113.065 ;
        RECT 115.705 112.555 116.385 113.125 ;
        RECT 118.895 112.555 119.575 113.125 ;
        RECT 50.500 104.060 106.660 105.560 ;
        RECT 128.875 88.885 157.175 89.515 ;
        RECT 156.545 8.265 157.175 88.885 ;
        RECT 156.560 1.000 157.160 8.265 ;
  END
END tt_um_mattvenn_r2r_dac
END LIBRARY

