module tt_um_prg_dup (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire \count[0] ;
 wire \count[1] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net3;
 wire net4;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire \out_count[0] ;
 wire \out_count[1] ;
 wire out_ready;
 wire \uut.R0[0] ;
 wire \uut.R0[1] ;
 wire \uut.R0[2] ;
 wire \uut.R0[3] ;
 wire \uut.R0[4] ;
 wire \uut.R0[5] ;
 wire \uut.R0[6] ;
 wire \uut.R0[7] ;
 wire \uut.R1[0] ;
 wire \uut.R1[1] ;
 wire \uut.R1[2] ;
 wire \uut.R1[3] ;
 wire \uut.R1[4] ;
 wire \uut.R1[5] ;
 wire \uut.R1[6] ;
 wire \uut.R1[7] ;
 wire \uut.in1[0] ;
 wire \uut.in1[1] ;
 wire \uut.in1[2] ;
 wire \uut.in1[3] ;
 wire \uut.in1[4] ;
 wire \uut.in1[5] ;
 wire \uut.in1[6] ;
 wire \uut.in1[7] ;
 wire \uut.in2[0] ;
 wire \uut.in2[1] ;
 wire \uut.in2[2] ;
 wire \uut.in2[3] ;
 wire \uut.in2[4] ;
 wire \uut.in2[5] ;
 wire \uut.in2[6] ;
 wire \uut.in2[7] ;
 wire \uut.in3[0] ;
 wire \uut.in3[1] ;
 wire \uut.in3[2] ;
 wire \uut.in3[3] ;
 wire \uut.in3[4] ;
 wire \uut.in3[5] ;
 wire \uut.in3[6] ;
 wire \uut.in3[7] ;
 wire \uut.mod_inv.inv_in1[0] ;
 wire \uut.mod_inv.inv_in1[1] ;
 wire \uut.mod_inv.inv_in1[2] ;
 wire \uut.mod_inv.inv_in1[3] ;
 wire \uut.mod_inv.inv_in2[0] ;
 wire \uut.mod_inv.inv_in2[1] ;
 wire \uut.mod_inv.inv_in2[2] ;
 wire \uut.mod_inv.inv_in2[3] ;
 wire \uut.mod_inv.inv_in3[0] ;
 wire \uut.mod_inv.inv_in3[1] ;
 wire \uut.mod_inv.inv_in3[2] ;
 wire \uut.mod_inv.inv_in3[3] ;
 wire \uut.mod_inv.inv_in4[0] ;
 wire \uut.mod_inv.inv_in4[1] ;
 wire \uut.mod_inv.inv_in4[2] ;
 wire \uut.mod_inv.inv_in4[3] ;
 wire \uut.mod_inv.inv_mod/_000_ ;
 wire \uut.mod_inv.inv_mod/_001_ ;
 wire \uut.mod_inv.inv_mod/_002_ ;
 wire \uut.mod_inv.inv_mod/_003_ ;
 wire \uut.mod_inv.inv_mod/_004_ ;
 wire \uut.mod_inv.inv_mod/_005_ ;
 wire \uut.mod_inv.inv_mod/_006_ ;
 wire \uut.mod_inv.inv_mod/_007_ ;
 wire \uut.mod_inv.inv_mod/_008_ ;
 wire \uut.mod_inv.inv_mod/_009_ ;
 wire \uut.mod_inv.inv_mod/_010_ ;
 wire \uut.mod_inv.inv_mod/_011_ ;
 wire \uut.mod_inv.inv_mod/_012_ ;
 wire \uut.mod_inv.inv_mod/_013_ ;
 wire \uut.mod_inv.inv_mod/_014_ ;
 wire \uut.mod_inv.inv_mod/_015_ ;
 wire \uut.mod_inv.inv_mod/_016_ ;
 wire \uut.mod_inv.inv_mod/_017_ ;
 wire \uut.mod_inv.inv_mod/_018_ ;
 wire \uut.mod_inv.inv_mod/_019_ ;
 wire \uut.mod_inv.inv_mod/_020_ ;
 wire \uut.mod_inv.inv_mod/_021_ ;
 wire \uut.mod_inv.inv_mod/_022_ ;
 wire \uut.mod_inv.inv_mod/_023_ ;
 wire \uut.mod_inv.inv_mod/_024_ ;
 wire \uut.mod_inv.inv_mod/_025_ ;
 wire \uut.mod_inv.inv_mod/_026_ ;
 wire \uut.mod_inv.inv_mod/_027_ ;
 wire \uut.mod_inv.inv_mod/_028_ ;
 wire \uut.mod_inv.inv_mod/_029_ ;
 wire \uut.mod_inv.inv_mod/_030_ ;
 wire \uut.mod_inv.inv_mod/_031_ ;
 wire \uut.mod_inv.inv_mod/_032_ ;
 wire \uut.mod_inv.inv_mod/_033_ ;
 wire \uut.mod_inv.inv_mod/_034_ ;
 wire \uut.mod_inv.inv_mod/_035_ ;
 wire \uut.mod_inv.inv_mod/_036_ ;
 wire \uut.mod_inv.inv_mod/_037_ ;
 wire \uut.mod_inv.inv_mod/_038_ ;
 wire \uut.mod_inv.inv_mod/_039_ ;
 wire \uut.mod_inv.inv_mod/_040_ ;
 wire \uut.mod_inv.inv_mod/_041_ ;
 wire \uut.mod_inv.inv_mod/_042_ ;
 wire \uut.mod_inv.inv_mod/_043_ ;
 wire \uut.mod_inv.inv_mod/_044_ ;
 wire \uut.mod_inv.inv_mod/_045_ ;
 wire \uut.mod_inv.inv_mod/_046_ ;
 wire \uut.mod_inv.inv_mod/_047_ ;
 wire \uut.mod_inv.inv_mod/_048_ ;
 wire \uut.mod_inv.inv_mod/_049_ ;
 wire \uut.mod_inv.inv_mod/_050_ ;
 wire \uut.mod_inv.inv_mod/_051_ ;
 wire \uut.mod_inv.inv_mod/_052_ ;
 wire \uut.mod_inv.inv_mod/_053_ ;
 wire \uut.mod_inv.inv_mod/_054_ ;
 wire \uut.mod_inv.inv_mod/_055_ ;
 wire \uut.mod_inv.inv_mod/_056_ ;
 wire \uut.mod_inv.inv_mod/_057_ ;
 wire \uut.mod_inv.inv_mod/_058_ ;
 wire \uut.mod_inv.inv_mod/_059_ ;
 wire \uut.mod_inv.inv_mod/_060_ ;
 wire \uut.mod_inv.inv_mod/_061_ ;
 wire \uut.mod_inv.inv_mod/_062_ ;
 wire \uut.mod_inv.inv_mod/_063_ ;
 wire \uut.mod_inv.inv_mod/_064_ ;
 wire \uut.mod_inv.inv_mod/_065_ ;
 wire \uut.mod_inv.inv_mod/_066_ ;
 wire \uut.mod_inv.inv_mod/_067_ ;
 wire \uut.mod_inv.inv_mod/_068_ ;
 wire \uut.mod_inv.inv_mod/_069_ ;
 wire \uut.mod_inv.inv_mod/_070_ ;
 wire \uut.mod_inv.inv_mod/_071_ ;
 wire \uut.mod_inv.inv_mod/_072_ ;
 wire \uut.mod_inv.inv_mod/_073_ ;
 wire \uut.mod_inv.inv_mod/_074_ ;
 wire \uut.mod_inv.inv_mod/_075_ ;
 wire \uut.mod_inv.inv_mod/_076_ ;
 wire \uut.mod_inv.inv_mod/_077_ ;
 wire \uut.mod_inv.inv_mod/_078_ ;
 wire \uut.mod_inv.inv_mod/_079_ ;
 wire \uut.mod_inv.inv_mod/_080_ ;
 wire \uut.mod_inv.inv_mod/_081_ ;
 wire \uut.mod_inv.inv_mod/_082_ ;
 wire \uut.mod_inv.inv_mod/_083_ ;
 wire \uut.mod_inv.inv_mod/_084_ ;
 wire \uut.mod_inv.inv_mod/_085_ ;
 wire \uut.mod_inv.inv_mod/_086_ ;
 wire \uut.mod_inv.inv_mod/_087_ ;
 wire \uut.mod_inv.inv_mod/_088_ ;
 wire \uut.mod_inv.inv_mod/_089_ ;
 wire \uut.mod_inv.inv_mod/_090_ ;
 wire \uut.mod_inv.inv_mod/_091_ ;
 wire \uut.mod_inv.inv_mod/_092_ ;
 wire \uut.mod_inv.inv_mod/_093_ ;
 wire \uut.mod_inv.inv_mod/_094_ ;
 wire \uut.mod_inv.inv_mod/_095_ ;
 wire \uut.mod_inv.inv_mod/_096_ ;
 wire \uut.mod_inv.inv_mod/_097_ ;
 wire \uut.mod_inv.inv_mod/_098_ ;
 wire \uut.mod_inv.inv_mod/_099_ ;
 wire \uut.mod_inv.inv_mod/_100_ ;
 wire \uut.mod_inv.inv_mod/_101_ ;
 wire \uut.mod_inv.inv_mod/_102_ ;
 wire \uut.mod_inv.inv_mod/_103_ ;
 wire \uut.mod_inv.inv_mod/_104_ ;
 wire \uut.mod_inv.inv_mod/_105_ ;
 wire \uut.mod_inv.inv_mod/_106_ ;
 wire \uut.mod_inv.inv_mod/_107_ ;
 wire \uut.mod_inv.inv_mod/_108_ ;
 wire \uut.mod_inv.inv_mod/_109_ ;
 wire \uut.mod_inv.inv_mod/_110_ ;
 wire \uut.mod_inv.inv_mod/_111_ ;
 wire \uut.mod_inv.inv_mod/_112_ ;
 wire \uut.mod_inv.inv_mod/_113_ ;
 wire \uut.mod_inv.inv_mod/_114_ ;
 wire \uut.mod_inv.inv_mod/_115_ ;
 wire \uut.mod_inv.inv_mod/_116_ ;
 wire \uut.mod_inv.inv_mod/_117_ ;
 wire \uut.mod_inv.inv_mod/_118_ ;
 wire \uut.mod_inv.inv_mod/_119_ ;
 wire \uut.mod_inv.inv_mod/_120_ ;
 wire \uut.mod_inv.inv_mod/_121_ ;
 wire \uut.mod_inv.inv_mod/_122_ ;
 wire \uut.mod_inv.inv_mod/_123_ ;
 wire \uut.mod_inv.inv_mod/_124_ ;
 wire \uut.mod_inv.inv_mod/_125_ ;
 wire \uut.mod_inv.inv_mod/_126_ ;
 wire \uut.mod_inv.inv_mod/_127_ ;
 wire \uut.mod_inv.inv_mod/_128_ ;
 wire \uut.mod_inv.inv_mod/_129_ ;
 wire \uut.mod_inv.inv_mod/_130_ ;
 wire \uut.mod_inv.inv_mod/_131_ ;
 wire \uut.mod_inv.inv_mod/_132_ ;
 wire \uut.mod_inv.inv_mod/_133_ ;
 wire \uut.mod_inv.inv_mod/_134_ ;
 wire \uut.mod_inv.inv_mod/_135_ ;
 wire \uut.mod_inv.inv_mod/_136_ ;
 wire \uut.mod_inv.inv_mod/_137_ ;
 wire \uut.mod_inv.inv_mod/_138_ ;
 wire \uut.mod_inv.inv_mod/_139_ ;
 wire \uut.mod_inv.inv_mod/_140_ ;
 wire \uut.mod_inv.inv_mod/_141_ ;
 wire \uut.mod_inv.inv_mod/_142_ ;
 wire \uut.mod_inv.inv_mod/_143_ ;
 wire \uut.mod_inv.inv_mod/_144_ ;
 wire \uut.mod_inv.inv_mod/_145_ ;
 wire \uut.mod_inv.inv_mod/_146_ ;
 wire \uut.mod_inv.inv_mod/_147_ ;
 wire \uut.mod_inv.inv_mod/_148_ ;
 wire \uut.mod_inv.inv_mod/_149_ ;
 wire \uut.mod_inv.inv_mod/_150_ ;
 wire \uut.mod_inv.inv_mod/_151_ ;
 wire \uut.mod_inv.inv_mod/_152_ ;
 wire \uut.mod_inv.inv_mod/_153_ ;
 wire \uut.mod_inv.inv_mod/_154_ ;
 wire \uut.mod_inv.inv_mod/_155_ ;
 wire \uut.mod_inv.inv_mod/_156_ ;
 wire \uut.mod_inv.inv_mod/_157_ ;
 wire \uut.mod_inv.inv_mod/_158_ ;
 wire \uut.mod_inv.inv_mod/_159_ ;
 wire \uut.mod_inv.inv_mod/_160_ ;
 wire \uut.mod_inv.inv_mod/_161_ ;
 wire \uut.mod_inv.inv_mod/_162_ ;
 wire \uut.mod_inv.inv_mod/_163_ ;
 wire \uut.mod_inv.inv_mod/_164_ ;
 wire \uut.mod_inv.inv_mod/_165_ ;
 wire \uut.mod_inv.inv_mod/_166_ ;
 wire \uut.mod_inv.inv_mod/_167_ ;
 wire \uut.mod_inv.inv_mod/_168_ ;
 wire \uut.mod_inv.inv_mod/_169_ ;
 wire \uut.mod_inv.inv_mod/_170_ ;
 wire \uut.mod_inv.inv_mod/_171_ ;
 wire \uut.mod_inv.inv_mod/_172_ ;
 wire \uut.mod_inv.inv_mod/_173_ ;
 wire \uut.mod_inv.inv_mod/_174_ ;
 wire \uut.mod_inv.inv_mod/_175_ ;
 wire \uut.mod_inv.inv_mod/_176_ ;
 wire \uut.mod_inv.inv_mod/_177_ ;
 wire \uut.mod_inv.inv_mod/_178_ ;
 wire \uut.mod_inv.inv_mod/_179_ ;
 wire \uut.mod_inv.inv_mod/_180_ ;
 wire \uut.mod_inv.inv_mod/_181_ ;
 wire \uut.mod_inv.inv_mod/_182_ ;
 wire \uut.mod_inv.inv_mod/_183_ ;
 wire \uut.mod_inv.inv_mod/_184_ ;
 wire \uut.mod_inv.inv_mod/_185_ ;
 wire \uut.mod_inv.inv_mod/_186_ ;
 wire \uut.mod_inv.inv_mod/_187_ ;
 wire \uut.mod_inv.inv_mod/_188_ ;
 wire \uut.mod_inv.inv_mod/_189_ ;
 wire \uut.mod_inv.inv_mod/_190_ ;
 wire \uut.mod_inv.inv_mod/_191_ ;
 wire \uut.mod_inv.inv_mod/_192_ ;
 wire \uut.mod_inv.inv_mod/_193_ ;
 wire \uut.mod_inv.inv_mod/_194_ ;
 wire \uut.mod_inv.inv_mod/_195_ ;
 wire \uut.mod_inv.inv_mod/_196_ ;
 wire \uut.mod_inv.inv_mod/_197_ ;
 wire \uut.mod_inv.inv_mod/_198_ ;
 wire \uut.mod_inv.inv_mod/_199_ ;
 wire \uut.mod_inv.inv_mod/_200_ ;
 wire \uut.mod_inv.inv_mod/_201_ ;
 wire \uut.mod_inv.inv_mod/_202_ ;
 wire \uut.mod_inv.inv_mod/_203_ ;
 wire \uut.mod_inv.inv_mod/_204_ ;
 wire \uut.mod_inv.inv_mod/_205_ ;
 wire \uut.mod_inv.inv_mod/_206_ ;
 wire \uut.mod_inv.inv_mod/_207_ ;
 wire \uut.mod_inv.inv_mod/_208_ ;
 wire \uut.mod_inv.inv_mod/_209_ ;
 wire \uut.mod_inv.inv_mod/_210_ ;
 wire \uut.mod_inv.inv_mod/_211_ ;
 wire \uut.mod_inv.inv_mod/_212_ ;
 wire \uut.mod_inv.inv_mod/_213_ ;
 wire \uut.mod_inv.inv_mod/_214_ ;
 wire \uut.mod_inv.inv_mod/_215_ ;
 wire \uut.mod_inv.inv_mod/_216_ ;
 wire \uut.mod_inv.inv_mod/_217_ ;
 wire \uut.mod_inv.inv_mod/_218_ ;
 wire \uut.mod_inv.inv_mod/_219_ ;
 wire \uut.mod_inv.inv_mod/_220_ ;
 wire \uut.mod_inv.inv_mod/_221_ ;
 wire \uut.mod_inv.inv_mod/_222_ ;
 wire \uut.mod_inv.inv_mod/_223_ ;
 wire \uut.mod_inv.inv_mod/_224_ ;
 wire \uut.mod_inv.inv_mod/_225_ ;
 wire \uut.mod_inv.inv_mod/_226_ ;
 wire \uut.mod_inv.inv_mod/_227_ ;
 wire \uut.mod_inv.inv_mod/_228_ ;
 wire \uut.mod_inv.inv_mod/_229_ ;
 wire \uut.mod_inv.inv_mod/_230_ ;
 wire \uut.mod_inv.inv_mod/_231_ ;
 wire \uut.mod_inv.inv_mod/_232_ ;
 wire \uut.mod_inv.inv_mod/_233_ ;
 wire \uut.mod_inv.inv_mod/_234_ ;
 wire \uut.mod_inv.inv_mod/_235_ ;
 wire \uut.mod_inv.inv_mod/_236_ ;
 wire \uut.mod_inv.inv_mod/_237_ ;
 wire \uut.mod_inv.inv_mod/_238_ ;
 wire \uut.mod_inv.inv_mod/_239_ ;
 wire \uut.mod_inv.inv_mod/_240_ ;
 wire \uut.mod_inv.inv_mod/_241_ ;
 wire \uut.mod_inv.inv_mod/_242_ ;
 wire \uut.mod_inv.inv_mod/_243_ ;
 wire \uut.mod_inv.inv_mod/_244_ ;
 wire \uut.mod_inv.inv_mod/_245_ ;
 wire \uut.mod_inv.inv_mod/_246_ ;
 wire \uut.mod_inv.inv_mod/_247_ ;
 wire \uut.mod_inv.inv_mod/_248_ ;
 wire \uut.mod_inv.inv_mod/_249_ ;
 wire \uut.mod_inv.inv_mod/_250_ ;
 wire \uut.mod_inv.inv_mod/_251_ ;
 wire \uut.mod_inv.inv_mod/_252_ ;
 wire \uut.mod_inv.inv_mod/_253_ ;
 wire \uut.mod_inv.inv_mod/_254_ ;
 wire \uut.mod_inv.inv_out1[0] ;
 wire \uut.mod_inv.inv_out1[1] ;
 wire \uut.mod_inv.inv_out1[2] ;
 wire \uut.mod_inv.inv_out1[3] ;
 wire \uut.mod_inv.inv_out1_reg[0] ;
 wire \uut.mod_inv.inv_out1_reg[1] ;
 wire \uut.mod_inv.inv_out1_reg[2] ;
 wire \uut.mod_inv.inv_out1_reg[3] ;
 wire \uut.mod_inv.inv_out2[0] ;
 wire \uut.mod_inv.inv_out2[1] ;
 wire \uut.mod_inv.inv_out2[2] ;
 wire \uut.mod_inv.inv_out2[3] ;
 wire \uut.mod_inv.inv_out2_xor[0] ;
 wire \uut.mod_inv.inv_out2_xor[1] ;
 wire \uut.mod_inv.inv_out2_xor[2] ;
 wire \uut.mod_inv.inv_out2_xor[3] ;
 wire \uut.mod_inv.inv_out3[0] ;
 wire \uut.mod_inv.inv_out3[1] ;
 wire \uut.mod_inv.inv_out3[2] ;
 wire \uut.mod_inv.inv_out3[3] ;
 wire \uut.mod_inv.inv_out3_xor[0] ;
 wire \uut.mod_inv.inv_out3_xor[1] ;
 wire \uut.mod_inv.inv_out3_xor[2] ;
 wire \uut.mod_inv.inv_out3_xor[3] ;
 wire \uut.mod_inv.inv_out4[0] ;
 wire \uut.mod_inv.inv_out4[1] ;
 wire \uut.mod_inv.inv_out4[2] ;
 wire \uut.mod_inv.inv_out4[3] ;
 wire \uut.mod_inv.inv_out4_reg[0] ;
 wire \uut.mod_inv.inv_out4_reg[1] ;
 wire \uut.mod_inv.inv_out4_reg[2] ;
 wire \uut.mod_inv.inv_out4_reg[3] ;
 wire \uut.mod_inv.mod_mul1/_000_ ;
 wire \uut.mod_inv.mod_mul1/_001_ ;
 wire \uut.mod_inv.mod_mul1/_002_ ;
 wire \uut.mod_inv.mod_mul1/_003_ ;
 wire \uut.mod_inv.mod_mul1/_004_ ;
 wire \uut.mod_inv.mod_mul1/_005_ ;
 wire \uut.mod_inv.mod_mul1/_006_ ;
 wire \uut.mod_inv.mod_mul1/_007_ ;
 wire \uut.mod_inv.mod_mul1/_008_ ;
 wire \uut.mod_inv.mod_mul1/_009_ ;
 wire \uut.mod_inv.mod_mul1/_010_ ;
 wire \uut.mod_inv.mod_mul1/_011_ ;
 wire \uut.mod_inv.mod_mul1/_012_ ;
 wire \uut.mod_inv.mod_mul1/_013_ ;
 wire \uut.mod_inv.mod_mul1/_014_ ;
 wire \uut.mod_inv.mod_mul1/_015_ ;
 wire \uut.mod_inv.mod_mul1/_016_ ;
 wire \uut.mod_inv.mod_mul1/_017_ ;
 wire \uut.mod_inv.mod_mul1/_018_ ;
 wire \uut.mod_inv.mod_mul1/_019_ ;
 wire \uut.mod_inv.mod_mul1/_020_ ;
 wire \uut.mod_inv.mod_mul1/_021_ ;
 wire \uut.mod_inv.mod_mul1/_022_ ;
 wire \uut.mod_inv.mod_mul1/_023_ ;
 wire \uut.mod_inv.mod_mul1/_024_ ;
 wire \uut.mod_inv.mod_mul1/_025_ ;
 wire \uut.mod_inv.mod_mul1/_026_ ;
 wire \uut.mod_inv.mod_mul1/_027_ ;
 wire \uut.mod_inv.mod_mul1/_028_ ;
 wire \uut.mod_inv.mod_mul1/_029_ ;
 wire \uut.mod_inv.mod_mul1/_030_ ;
 wire \uut.mod_inv.mod_mul1/_031_ ;
 wire \uut.mod_inv.mod_mul1/_032_ ;
 wire \uut.mod_inv.mod_mul1/_033_ ;
 wire \uut.mod_inv.mod_mul1/_034_ ;
 wire \uut.mod_inv.mod_mul1/_035_ ;
 wire \uut.mod_inv.mod_mul1/_036_ ;
 wire \uut.mod_inv.mod_mul1/_037_ ;
 wire \uut.mod_inv.mod_mul1/_038_ ;
 wire \uut.mod_inv.mod_mul1/_039_ ;
 wire \uut.mod_inv.mod_mul1/_040_ ;
 wire \uut.mod_inv.mod_mul1/_041_ ;
 wire \uut.mod_inv.mod_mul1/_042_ ;
 wire \uut.mod_inv.mod_mul1/_043_ ;
 wire \uut.mod_inv.mod_mul1/_044_ ;
 wire \uut.mod_inv.mod_mul1/_045_ ;
 wire \uut.mod_inv.mod_mul1/_046_ ;
 wire \uut.mod_inv.mod_mul1/_047_ ;
 wire \uut.mod_inv.mod_mul1/_048_ ;
 wire \uut.mod_inv.mod_mul1/_049_ ;
 wire \uut.mod_inv.mod_mul1/_050_ ;
 wire \uut.mod_inv.mod_mul1/_051_ ;
 wire \uut.mod_inv.mod_mul1/_052_ ;
 wire \uut.mod_inv.mod_mul1/_053_ ;
 wire \uut.mod_inv.mod_mul1/_054_ ;
 wire \uut.mod_inv.mod_mul1/_055_ ;
 wire \uut.mod_inv.mod_mul1/_056_ ;
 wire \uut.mod_inv.mod_mul1/_057_ ;
 wire \uut.mod_inv.mod_mul1/_058_ ;
 wire \uut.mod_inv.mod_mul1/_059_ ;
 wire \uut.mod_inv.mod_mul1/_060_ ;
 wire \uut.mod_inv.mod_mul1/_061_ ;
 wire \uut.mod_inv.mod_mul1/_062_ ;
 wire \uut.mod_inv.mod_mul1/_063_ ;
 wire \uut.mod_inv.mod_mul1/_064_ ;
 wire \uut.mod_inv.mod_mul1/_065_ ;
 wire \uut.mod_inv.mod_mul1/_066_ ;
 wire \uut.mod_inv.mod_mul1/_067_ ;
 wire \uut.mod_inv.mod_mul1/_068_ ;
 wire \uut.mod_inv.mod_mul1/_069_ ;
 wire \uut.mod_inv.mod_mul1/_070_ ;
 wire \uut.mod_inv.mod_mul1/_071_ ;
 wire \uut.mod_inv.mod_mul1/_072_ ;
 wire \uut.mod_inv.mod_mul1/_073_ ;
 wire \uut.mod_inv.mod_mul1/_074_ ;
 wire \uut.mod_inv.mod_mul1/_075_ ;
 wire \uut.mod_inv.mod_mul1/_076_ ;
 wire \uut.mod_inv.mod_mul1/_077_ ;
 wire \uut.mod_inv.mod_mul1/_078_ ;
 wire \uut.mod_inv.mod_mul1/_079_ ;
 wire \uut.mod_inv.mod_mul1/_080_ ;
 wire \uut.mod_inv.mod_mul1/_081_ ;
 wire \uut.mod_inv.mod_mul1/_082_ ;
 wire \uut.mod_inv.mod_mul1/_083_ ;
 wire \uut.mod_inv.mod_mul1/_084_ ;
 wire \uut.mod_inv.mod_mul1/_085_ ;
 wire \uut.mod_inv.mod_mul1/_086_ ;
 wire \uut.mod_inv.mod_mul1/_087_ ;
 wire \uut.mod_inv.mod_mul1/_088_ ;
 wire \uut.mod_inv.mod_mul1/_089_ ;
 wire \uut.mod_inv.mod_mul1/_090_ ;
 wire \uut.mod_inv.mod_mul1/_091_ ;
 wire \uut.mod_inv.mod_mul1/_092_ ;
 wire \uut.mod_inv.mod_mul1/_093_ ;
 wire \uut.mod_inv.mod_mul1/_094_ ;
 wire \uut.mod_inv.mod_mul1/_095_ ;
 wire \uut.mod_inv.mod_mul1/_096_ ;
 wire \uut.mod_inv.mod_mul1/_097_ ;
 wire \uut.mod_inv.mod_mul1/_098_ ;
 wire \uut.mod_inv.mod_mul1/_099_ ;
 wire \uut.mod_inv.mod_mul1/_100_ ;
 wire \uut.mod_inv.mod_mul1/_101_ ;
 wire \uut.mod_inv.mod_mul1/_102_ ;
 wire \uut.mod_inv.mod_mul1/_103_ ;
 wire \uut.mod_inv.mod_mul1/_104_ ;
 wire \uut.mod_inv.mod_mul1/_105_ ;
 wire \uut.mod_inv.mod_mul1/_106_ ;
 wire \uut.mod_inv.mod_mul1/_107_ ;
 wire \uut.mod_inv.mod_mul1/_108_ ;
 wire \uut.mod_inv.mod_mul1/_109_ ;
 wire \uut.mod_inv.mod_mul1/_110_ ;
 wire \uut.mod_inv.mod_mul1/_111_ ;
 wire \uut.mod_inv.mod_mul1/_112_ ;
 wire \uut.mod_inv.mod_mul1/_113_ ;
 wire \uut.mod_inv.mod_mul1/_114_ ;
 wire \uut.mod_inv.mod_mul1/_115_ ;
 wire \uut.mod_inv.mod_mul1/_116_ ;
 wire \uut.mod_inv.mod_mul1/_117_ ;
 wire \uut.mod_inv.mod_mul1/_118_ ;
 wire \uut.mod_inv.mod_mul1/_119_ ;
 wire \uut.mod_inv.mod_mul1/_120_ ;
 wire \uut.mod_inv.mod_mul1/_121_ ;
 wire \uut.mod_inv.mod_mul1/_122_ ;
 wire \uut.mod_inv.mod_mul1/_123_ ;
 wire \uut.mod_inv.mod_mul1/_124_ ;
 wire \uut.mod_inv.mod_mul1/_125_ ;
 wire \uut.mod_inv.mod_mul1/_126_ ;
 wire \uut.mod_inv.mod_mul1/_127_ ;
 wire \uut.mod_inv.mod_mul1/_128_ ;
 wire \uut.mod_inv.mod_mul1/_129_ ;
 wire \uut.mod_inv.mod_mul1/_130_ ;
 wire \uut.mod_inv.mod_mul1/_131_ ;
 wire \uut.mod_inv.mod_mul1/_132_ ;
 wire \uut.mod_inv.mod_mul1/_133_ ;
 wire \uut.mod_inv.mod_mul1/_134_ ;
 wire \uut.mod_inv.mod_mul1/_135_ ;
 wire \uut.mod_inv.mod_mul1/_136_ ;
 wire \uut.mod_inv.mod_mul1/_137_ ;
 wire \uut.mod_inv.mod_mul1/_138_ ;
 wire \uut.mod_inv.mod_mul1/_139_ ;
 wire \uut.mod_inv.mod_mul1/_140_ ;
 wire \uut.mod_inv.mod_mul1/_141_ ;
 wire \uut.mod_inv.mod_mul1/_142_ ;
 wire \uut.mod_inv.mod_mul1/_143_ ;
 wire \uut.mod_inv.mod_mul1/_144_ ;
 wire \uut.mod_inv.mod_mul1/_145_ ;
 wire \uut.mod_inv.mod_mul1/_146_ ;
 wire \uut.mod_inv.mod_mul1/_147_ ;
 wire \uut.mod_inv.mod_mul1/_148_ ;
 wire \uut.mod_inv.mod_mul1/_149_ ;
 wire \uut.mod_inv.mod_mul1/_150_ ;
 wire \uut.mod_inv.mod_mul1/_151_ ;
 wire \uut.mod_inv.mod_mul1/_152_ ;
 wire \uut.mod_inv.mod_mul1/_153_ ;
 wire \uut.mod_inv.mod_mul1/_154_ ;
 wire \uut.mod_inv.mod_mul1/_155_ ;
 wire \uut.mod_inv.mod_mul1/_156_ ;
 wire \uut.mod_inv.mod_mul1/_157_ ;
 wire \uut.mod_inv.mod_mul1/_158_ ;
 wire \uut.mod_inv.mod_mul1/_159_ ;
 wire \uut.mod_inv.mod_mul1/_160_ ;
 wire \uut.mod_inv.mod_mul1/_161_ ;
 wire \uut.mod_inv.mod_mul1/_162_ ;
 wire \uut.mod_inv.mod_mul1/_163_ ;
 wire \uut.mod_inv.mod_mul1/_164_ ;
 wire \uut.mod_inv.mod_mul1/_165_ ;
 wire \uut.mod_inv.mod_mul1/_166_ ;
 wire \uut.mod_inv.mod_mul1/_167_ ;
 wire \uut.mod_inv.mod_mul1/_168_ ;
 wire \uut.mod_inv.mod_mul1/_169_ ;
 wire \uut.mod_inv.mod_mul1/_170_ ;
 wire \uut.mod_inv.mod_mul1/_171_ ;
 wire \uut.mod_inv.mod_mul1/_172_ ;
 wire \uut.mod_inv.mod_mul1/_173_ ;
 wire \uut.mod_inv.mod_mul1/_174_ ;
 wire \uut.mod_inv.mod_mul1/_175_ ;
 wire \uut.mod_inv.mod_mul1/_176_ ;
 wire \uut.mod_inv.mod_mul1/_177_ ;
 wire \uut.mod_inv.mod_mul1/_178_ ;
 wire \uut.mod_inv.mod_mul1/_179_ ;
 wire \uut.mod_inv.mod_mul1/_180_ ;
 wire \uut.mod_inv.mod_mul1/_181_ ;
 wire \uut.mod_inv.mod_mul1/_182_ ;
 wire \uut.mod_inv.mod_mul1/_183_ ;
 wire \uut.mod_inv.mod_mul1/_184_ ;
 wire \uut.mod_inv.mod_mul1/_185_ ;
 wire \uut.mod_inv.mod_mul1/_186_ ;
 wire \uut.mod_inv.mod_mul1/_187_ ;
 wire \uut.mod_inv.mod_mul1/_188_ ;
 wire \uut.mod_inv.mod_mul1/_189_ ;
 wire \uut.mod_inv.mod_mul1/_190_ ;
 wire \uut.mod_inv.mod_mul1/_191_ ;
 wire \uut.mod_inv.mod_mul1/_192_ ;
 wire \uut.mod_inv.mod_mul1/_193_ ;
 wire \uut.mod_inv.mod_mul1/_194_ ;
 wire \uut.mod_inv.mod_mul1/_195_ ;
 wire \uut.mod_inv.mod_mul1/_196_ ;
 wire \uut.mod_inv.mod_mul1/_197_ ;
 wire \uut.mod_inv.mod_mul1/_198_ ;
 wire \uut.mod_inv.mod_mul1/_199_ ;
 wire \uut.mod_inv.mod_mul1/_200_ ;
 wire \uut.mod_inv.mod_mul1/_201_ ;
 wire \uut.mod_inv.mod_mul1/_202_ ;
 wire \uut.mod_inv.mod_mul1/_203_ ;
 wire \uut.mod_inv.mod_mul1/_204_ ;
 wire \uut.mod_inv.mod_mul1/_205_ ;
 wire \uut.mod_inv.mod_mul1/_206_ ;
 wire \uut.mod_inv.mod_mul1/_207_ ;
 wire \uut.mod_inv.mod_mul1/_208_ ;
 wire \uut.mod_inv.mod_mul1/_209_ ;
 wire \uut.mod_inv.mod_mul1/_210_ ;
 wire \uut.mod_inv.mod_mul1/_211_ ;
 wire \uut.mod_inv.mod_mul1/_212_ ;
 wire \uut.mod_inv.mod_mul1/_213_ ;
 wire \uut.mod_inv.mod_mul1/_214_ ;
 wire \uut.mod_inv.mod_mul1/_215_ ;
 wire \uut.mod_inv.mod_mul1/_216_ ;
 wire \uut.mod_inv.mod_mul1/_217_ ;
 wire \uut.mod_inv.mod_mul1/_218_ ;
 wire \uut.mod_inv.mod_mul1/_219_ ;
 wire \uut.mod_inv.mod_mul1/_220_ ;
 wire \uut.mod_inv.mod_mul1_out1[0] ;
 wire \uut.mod_inv.mod_mul1_out1[1] ;
 wire \uut.mod_inv.mod_mul1_out1[2] ;
 wire \uut.mod_inv.mod_mul1_out1[3] ;
 wire \uut.mod_inv.mod_mul1_out1_reg[0] ;
 wire \uut.mod_inv.mod_mul1_out1_reg[1] ;
 wire \uut.mod_inv.mod_mul1_out1_reg[2] ;
 wire \uut.mod_inv.mod_mul1_out1_reg[3] ;
 wire \uut.mod_inv.mod_mul1_out2[0] ;
 wire \uut.mod_inv.mod_mul1_out2[1] ;
 wire \uut.mod_inv.mod_mul1_out2[2] ;
 wire \uut.mod_inv.mod_mul1_out2[3] ;
 wire \uut.mod_inv.mod_mul1_out2_xor[0] ;
 wire \uut.mod_inv.mod_mul1_out2_xor[1] ;
 wire \uut.mod_inv.mod_mul1_out2_xor[2] ;
 wire \uut.mod_inv.mod_mul1_out2_xor[3] ;
 wire \uut.mod_inv.mod_mul1_out3[0] ;
 wire \uut.mod_inv.mod_mul1_out3[1] ;
 wire \uut.mod_inv.mod_mul1_out3[2] ;
 wire \uut.mod_inv.mod_mul1_out3[3] ;
 wire \uut.mod_inv.mod_mul2/_000_ ;
 wire \uut.mod_inv.mod_mul2/_001_ ;
 wire \uut.mod_inv.mod_mul2/_002_ ;
 wire \uut.mod_inv.mod_mul2/_003_ ;
 wire \uut.mod_inv.mod_mul2/_004_ ;
 wire \uut.mod_inv.mod_mul2/_005_ ;
 wire \uut.mod_inv.mod_mul2/_006_ ;
 wire \uut.mod_inv.mod_mul2/_007_ ;
 wire \uut.mod_inv.mod_mul2/_008_ ;
 wire \uut.mod_inv.mod_mul2/_009_ ;
 wire \uut.mod_inv.mod_mul2/_010_ ;
 wire \uut.mod_inv.mod_mul2/_011_ ;
 wire \uut.mod_inv.mod_mul2/_012_ ;
 wire \uut.mod_inv.mod_mul2/_013_ ;
 wire \uut.mod_inv.mod_mul2/_014_ ;
 wire \uut.mod_inv.mod_mul2/_015_ ;
 wire \uut.mod_inv.mod_mul2/_016_ ;
 wire \uut.mod_inv.mod_mul2/_017_ ;
 wire \uut.mod_inv.mod_mul2/_018_ ;
 wire \uut.mod_inv.mod_mul2/_019_ ;
 wire \uut.mod_inv.mod_mul2/_020_ ;
 wire \uut.mod_inv.mod_mul2/_021_ ;
 wire \uut.mod_inv.mod_mul2/_022_ ;
 wire \uut.mod_inv.mod_mul2/_023_ ;
 wire \uut.mod_inv.mod_mul2/_024_ ;
 wire \uut.mod_inv.mod_mul2/_025_ ;
 wire \uut.mod_inv.mod_mul2/_026_ ;
 wire \uut.mod_inv.mod_mul2/_027_ ;
 wire \uut.mod_inv.mod_mul2/_028_ ;
 wire \uut.mod_inv.mod_mul2/_029_ ;
 wire \uut.mod_inv.mod_mul2/_030_ ;
 wire \uut.mod_inv.mod_mul2/_031_ ;
 wire \uut.mod_inv.mod_mul2/_032_ ;
 wire \uut.mod_inv.mod_mul2/_033_ ;
 wire \uut.mod_inv.mod_mul2/_034_ ;
 wire \uut.mod_inv.mod_mul2/_035_ ;
 wire \uut.mod_inv.mod_mul2/_036_ ;
 wire \uut.mod_inv.mod_mul2/_037_ ;
 wire \uut.mod_inv.mod_mul2/_038_ ;
 wire \uut.mod_inv.mod_mul2/_039_ ;
 wire \uut.mod_inv.mod_mul2/_040_ ;
 wire \uut.mod_inv.mod_mul2/_041_ ;
 wire \uut.mod_inv.mod_mul2/_042_ ;
 wire \uut.mod_inv.mod_mul2/_043_ ;
 wire \uut.mod_inv.mod_mul2/_044_ ;
 wire \uut.mod_inv.mod_mul2/_045_ ;
 wire \uut.mod_inv.mod_mul2/_046_ ;
 wire \uut.mod_inv.mod_mul2/_047_ ;
 wire \uut.mod_inv.mod_mul2/_048_ ;
 wire \uut.mod_inv.mod_mul2/_049_ ;
 wire \uut.mod_inv.mod_mul2/_050_ ;
 wire \uut.mod_inv.mod_mul2/_051_ ;
 wire \uut.mod_inv.mod_mul2/_052_ ;
 wire \uut.mod_inv.mod_mul2/_053_ ;
 wire \uut.mod_inv.mod_mul2/_054_ ;
 wire \uut.mod_inv.mod_mul2/_055_ ;
 wire \uut.mod_inv.mod_mul2/_056_ ;
 wire \uut.mod_inv.mod_mul2/_057_ ;
 wire \uut.mod_inv.mod_mul2/_058_ ;
 wire \uut.mod_inv.mod_mul2/_059_ ;
 wire \uut.mod_inv.mod_mul2/_060_ ;
 wire \uut.mod_inv.mod_mul2/_061_ ;
 wire \uut.mod_inv.mod_mul2/_062_ ;
 wire \uut.mod_inv.mod_mul2/_063_ ;
 wire \uut.mod_inv.mod_mul2/_064_ ;
 wire \uut.mod_inv.mod_mul2/_065_ ;
 wire \uut.mod_inv.mod_mul2/_066_ ;
 wire \uut.mod_inv.mod_mul2/_067_ ;
 wire \uut.mod_inv.mod_mul2/_068_ ;
 wire \uut.mod_inv.mod_mul2/_069_ ;
 wire \uut.mod_inv.mod_mul2/_070_ ;
 wire \uut.mod_inv.mod_mul2/_071_ ;
 wire \uut.mod_inv.mod_mul2/_072_ ;
 wire \uut.mod_inv.mod_mul2/_073_ ;
 wire \uut.mod_inv.mod_mul2/_074_ ;
 wire \uut.mod_inv.mod_mul2/_075_ ;
 wire \uut.mod_inv.mod_mul2/_076_ ;
 wire \uut.mod_inv.mod_mul2/_077_ ;
 wire \uut.mod_inv.mod_mul2/_078_ ;
 wire \uut.mod_inv.mod_mul2/_079_ ;
 wire \uut.mod_inv.mod_mul2/_080_ ;
 wire \uut.mod_inv.mod_mul2/_081_ ;
 wire \uut.mod_inv.mod_mul2/_082_ ;
 wire \uut.mod_inv.mod_mul2/_083_ ;
 wire \uut.mod_inv.mod_mul2/_084_ ;
 wire \uut.mod_inv.mod_mul2/_085_ ;
 wire \uut.mod_inv.mod_mul2/_086_ ;
 wire \uut.mod_inv.mod_mul2/_087_ ;
 wire \uut.mod_inv.mod_mul2/_088_ ;
 wire \uut.mod_inv.mod_mul2/_089_ ;
 wire \uut.mod_inv.mod_mul2/_090_ ;
 wire \uut.mod_inv.mod_mul2/_091_ ;
 wire \uut.mod_inv.mod_mul2/_092_ ;
 wire \uut.mod_inv.mod_mul2/_093_ ;
 wire \uut.mod_inv.mod_mul2/_094_ ;
 wire \uut.mod_inv.mod_mul2/_095_ ;
 wire \uut.mod_inv.mod_mul2/_096_ ;
 wire \uut.mod_inv.mod_mul2/_097_ ;
 wire \uut.mod_inv.mod_mul2/_098_ ;
 wire \uut.mod_inv.mod_mul2/_099_ ;
 wire \uut.mod_inv.mod_mul2/_100_ ;
 wire \uut.mod_inv.mod_mul2/_101_ ;
 wire \uut.mod_inv.mod_mul2/_102_ ;
 wire \uut.mod_inv.mod_mul2/_103_ ;
 wire \uut.mod_inv.mod_mul2/_104_ ;
 wire \uut.mod_inv.mod_mul2/_105_ ;
 wire \uut.mod_inv.mod_mul2/_106_ ;
 wire \uut.mod_inv.mod_mul2/_107_ ;
 wire \uut.mod_inv.mod_mul2/_108_ ;
 wire \uut.mod_inv.mod_mul2/_109_ ;
 wire \uut.mod_inv.mod_mul2/_110_ ;
 wire \uut.mod_inv.mod_mul2/_111_ ;
 wire \uut.mod_inv.mod_mul2/_112_ ;
 wire \uut.mod_inv.mod_mul2/_113_ ;
 wire \uut.mod_inv.mod_mul2/_114_ ;
 wire \uut.mod_inv.mod_mul2/_115_ ;
 wire \uut.mod_inv.mod_mul2/_116_ ;
 wire \uut.mod_inv.mod_mul2/_117_ ;
 wire \uut.mod_inv.mod_mul2/_118_ ;
 wire \uut.mod_inv.mod_mul2/_119_ ;
 wire \uut.mod_inv.mod_mul2/_120_ ;
 wire \uut.mod_inv.mod_mul2/_121_ ;
 wire \uut.mod_inv.mod_mul2/_122_ ;
 wire \uut.mod_inv.mod_mul2/_123_ ;
 wire \uut.mod_inv.mod_mul2/_124_ ;
 wire \uut.mod_inv.mod_mul2/_125_ ;
 wire \uut.mod_inv.mod_mul2/_126_ ;
 wire \uut.mod_inv.mod_mul2/_127_ ;
 wire \uut.mod_inv.mod_mul2/_128_ ;
 wire \uut.mod_inv.mod_mul2/_129_ ;
 wire \uut.mod_inv.mod_mul2/_130_ ;
 wire \uut.mod_inv.mod_mul2/_131_ ;
 wire \uut.mod_inv.mod_mul2/_132_ ;
 wire \uut.mod_inv.mod_mul2/_133_ ;
 wire \uut.mod_inv.mod_mul2/_134_ ;
 wire \uut.mod_inv.mod_mul2/_135_ ;
 wire \uut.mod_inv.mod_mul2/_136_ ;
 wire \uut.mod_inv.mod_mul2/_137_ ;
 wire \uut.mod_inv.mod_mul2/_138_ ;
 wire \uut.mod_inv.mod_mul2/_139_ ;
 wire \uut.mod_inv.mod_mul2/_140_ ;
 wire \uut.mod_inv.mod_mul2/_141_ ;
 wire \uut.mod_inv.mod_mul2/_142_ ;
 wire \uut.mod_inv.mod_mul2/_143_ ;
 wire \uut.mod_inv.mod_mul2/_144_ ;
 wire \uut.mod_inv.mod_mul2/_145_ ;
 wire \uut.mod_inv.mod_mul2/_146_ ;
 wire \uut.mod_inv.mod_mul2/_147_ ;
 wire \uut.mod_inv.mod_mul2/_148_ ;
 wire \uut.mod_inv.mod_mul2/_149_ ;
 wire \uut.mod_inv.mod_mul2/_150_ ;
 wire \uut.mod_inv.mod_mul2/_151_ ;
 wire \uut.mod_inv.mod_mul2/_152_ ;
 wire \uut.mod_inv.mod_mul2/_153_ ;
 wire \uut.mod_inv.mod_mul2/_154_ ;
 wire \uut.mod_inv.mod_mul2/_155_ ;
 wire \uut.mod_inv.mod_mul2/_156_ ;
 wire \uut.mod_inv.mod_mul2/_157_ ;
 wire \uut.mod_inv.mod_mul2/_158_ ;
 wire \uut.mod_inv.mod_mul2/_159_ ;
 wire \uut.mod_inv.mod_mul2/_160_ ;
 wire \uut.mod_inv.mod_mul2/_161_ ;
 wire \uut.mod_inv.mod_mul2/_162_ ;
 wire \uut.mod_inv.mod_mul2/_163_ ;
 wire \uut.mod_inv.mod_mul2/_164_ ;
 wire \uut.mod_inv.mod_mul2/_165_ ;
 wire \uut.mod_inv.mod_mul2/_166_ ;
 wire \uut.mod_inv.mod_mul2/_167_ ;
 wire \uut.mod_inv.mod_mul2/_168_ ;
 wire \uut.mod_inv.mod_mul2/_169_ ;
 wire \uut.mod_inv.mod_mul2/_170_ ;
 wire \uut.mod_inv.mod_mul2/_171_ ;
 wire \uut.mod_inv.mod_mul2/_172_ ;
 wire \uut.mod_inv.mod_mul2/_173_ ;
 wire \uut.mod_inv.mod_mul2/_174_ ;
 wire \uut.mod_inv.mod_mul2/_175_ ;
 wire \uut.mod_inv.mod_mul2/_176_ ;
 wire \uut.mod_inv.mod_mul2/_177_ ;
 wire \uut.mod_inv.mod_mul2/_178_ ;
 wire \uut.mod_inv.mod_mul2/_179_ ;
 wire \uut.mod_inv.mod_mul2/_180_ ;
 wire \uut.mod_inv.mod_mul2/_181_ ;
 wire \uut.mod_inv.mod_mul2/_182_ ;
 wire \uut.mod_inv.mod_mul2/_183_ ;
 wire \uut.mod_inv.mod_mul2/_184_ ;
 wire \uut.mod_inv.mod_mul2/_185_ ;
 wire \uut.mod_inv.mod_mul2/_186_ ;
 wire \uut.mod_inv.mod_mul2/_187_ ;
 wire \uut.mod_inv.mod_mul2/_188_ ;
 wire \uut.mod_inv.mod_mul2/_189_ ;
 wire \uut.mod_inv.mod_mul2/_190_ ;
 wire \uut.mod_inv.mod_mul2/_191_ ;
 wire \uut.mod_inv.mod_mul2/_192_ ;
 wire \uut.mod_inv.mod_mul2/_193_ ;
 wire \uut.mod_inv.mod_mul2/_194_ ;
 wire \uut.mod_inv.mod_mul2/_195_ ;
 wire \uut.mod_inv.mod_mul2/_196_ ;
 wire \uut.mod_inv.mod_mul2/_197_ ;
 wire \uut.mod_inv.mod_mul2/_198_ ;
 wire \uut.mod_inv.mod_mul2/_199_ ;
 wire \uut.mod_inv.mod_mul2/_200_ ;
 wire \uut.mod_inv.mod_mul2/_201_ ;
 wire \uut.mod_inv.mod_mul2/_202_ ;
 wire \uut.mod_inv.mod_mul2/_203_ ;
 wire \uut.mod_inv.mod_mul2/_204_ ;
 wire \uut.mod_inv.mod_mul2/_205_ ;
 wire \uut.mod_inv.mod_mul2/_206_ ;
 wire \uut.mod_inv.mod_mul2/_207_ ;
 wire \uut.mod_inv.mod_mul2/_208_ ;
 wire \uut.mod_inv.mod_mul2/_209_ ;
 wire \uut.mod_inv.mod_mul2/_210_ ;
 wire \uut.mod_inv.mod_mul2/_211_ ;
 wire \uut.mod_inv.mod_mul2/_212_ ;
 wire \uut.mod_inv.mod_mul2/_213_ ;
 wire \uut.mod_inv.mod_mul2/_214_ ;
 wire \uut.mod_inv.mod_mul2/_215_ ;
 wire \uut.mod_inv.mod_mul2/_216_ ;
 wire \uut.mod_inv.mod_mul2/_217_ ;
 wire \uut.mod_inv.mod_mul2/_218_ ;
 wire \uut.mod_inv.mod_mul2/_219_ ;
 wire \uut.mod_inv.mod_mul2/_220_ ;
 wire \uut.mod_inv.mod_mul2_out1[0] ;
 wire \uut.mod_inv.mod_mul2_out1[1] ;
 wire \uut.mod_inv.mod_mul2_out1[2] ;
 wire \uut.mod_inv.mod_mul2_out1[3] ;
 wire \uut.mod_inv.mod_mul2_out2[0] ;
 wire \uut.mod_inv.mod_mul2_out2[1] ;
 wire \uut.mod_inv.mod_mul2_out2[2] ;
 wire \uut.mod_inv.mod_mul2_out2[3] ;
 wire \uut.mod_inv.mod_mul2_out3[0] ;
 wire \uut.mod_inv.mod_mul2_out3[1] ;
 wire \uut.mod_inv.mod_mul2_out3[2] ;
 wire \uut.mod_inv.mod_mul2_out3[3] ;
 wire \uut.mod_inv.mod_mul3/_000_ ;
 wire \uut.mod_inv.mod_mul3/_001_ ;
 wire \uut.mod_inv.mod_mul3/_002_ ;
 wire \uut.mod_inv.mod_mul3/_003_ ;
 wire \uut.mod_inv.mod_mul3/_004_ ;
 wire \uut.mod_inv.mod_mul3/_005_ ;
 wire \uut.mod_inv.mod_mul3/_006_ ;
 wire \uut.mod_inv.mod_mul3/_007_ ;
 wire \uut.mod_inv.mod_mul3/_008_ ;
 wire \uut.mod_inv.mod_mul3/_009_ ;
 wire \uut.mod_inv.mod_mul3/_010_ ;
 wire \uut.mod_inv.mod_mul3/_011_ ;
 wire \uut.mod_inv.mod_mul3/_012_ ;
 wire \uut.mod_inv.mod_mul3/_013_ ;
 wire \uut.mod_inv.mod_mul3/_014_ ;
 wire \uut.mod_inv.mod_mul3/_015_ ;
 wire \uut.mod_inv.mod_mul3/_016_ ;
 wire \uut.mod_inv.mod_mul3/_017_ ;
 wire \uut.mod_inv.mod_mul3/_018_ ;
 wire \uut.mod_inv.mod_mul3/_019_ ;
 wire \uut.mod_inv.mod_mul3/_020_ ;
 wire \uut.mod_inv.mod_mul3/_021_ ;
 wire \uut.mod_inv.mod_mul3/_022_ ;
 wire \uut.mod_inv.mod_mul3/_023_ ;
 wire \uut.mod_inv.mod_mul3/_024_ ;
 wire \uut.mod_inv.mod_mul3/_025_ ;
 wire \uut.mod_inv.mod_mul3/_026_ ;
 wire \uut.mod_inv.mod_mul3/_027_ ;
 wire \uut.mod_inv.mod_mul3/_028_ ;
 wire \uut.mod_inv.mod_mul3/_029_ ;
 wire \uut.mod_inv.mod_mul3/_030_ ;
 wire \uut.mod_inv.mod_mul3/_031_ ;
 wire \uut.mod_inv.mod_mul3/_032_ ;
 wire \uut.mod_inv.mod_mul3/_033_ ;
 wire \uut.mod_inv.mod_mul3/_034_ ;
 wire \uut.mod_inv.mod_mul3/_035_ ;
 wire \uut.mod_inv.mod_mul3/_036_ ;
 wire \uut.mod_inv.mod_mul3/_037_ ;
 wire \uut.mod_inv.mod_mul3/_038_ ;
 wire \uut.mod_inv.mod_mul3/_039_ ;
 wire \uut.mod_inv.mod_mul3/_040_ ;
 wire \uut.mod_inv.mod_mul3/_041_ ;
 wire \uut.mod_inv.mod_mul3/_042_ ;
 wire \uut.mod_inv.mod_mul3/_043_ ;
 wire \uut.mod_inv.mod_mul3/_044_ ;
 wire \uut.mod_inv.mod_mul3/_045_ ;
 wire \uut.mod_inv.mod_mul3/_046_ ;
 wire \uut.mod_inv.mod_mul3/_047_ ;
 wire \uut.mod_inv.mod_mul3/_048_ ;
 wire \uut.mod_inv.mod_mul3/_049_ ;
 wire \uut.mod_inv.mod_mul3/_050_ ;
 wire \uut.mod_inv.mod_mul3/_051_ ;
 wire \uut.mod_inv.mod_mul3/_052_ ;
 wire \uut.mod_inv.mod_mul3/_053_ ;
 wire \uut.mod_inv.mod_mul3/_054_ ;
 wire \uut.mod_inv.mod_mul3/_055_ ;
 wire \uut.mod_inv.mod_mul3/_056_ ;
 wire \uut.mod_inv.mod_mul3/_057_ ;
 wire \uut.mod_inv.mod_mul3/_058_ ;
 wire \uut.mod_inv.mod_mul3/_059_ ;
 wire \uut.mod_inv.mod_mul3/_060_ ;
 wire \uut.mod_inv.mod_mul3/_061_ ;
 wire \uut.mod_inv.mod_mul3/_062_ ;
 wire \uut.mod_inv.mod_mul3/_063_ ;
 wire \uut.mod_inv.mod_mul3/_064_ ;
 wire \uut.mod_inv.mod_mul3/_065_ ;
 wire \uut.mod_inv.mod_mul3/_066_ ;
 wire \uut.mod_inv.mod_mul3/_067_ ;
 wire \uut.mod_inv.mod_mul3/_068_ ;
 wire \uut.mod_inv.mod_mul3/_069_ ;
 wire \uut.mod_inv.mod_mul3/_070_ ;
 wire \uut.mod_inv.mod_mul3/_071_ ;
 wire \uut.mod_inv.mod_mul3/_072_ ;
 wire \uut.mod_inv.mod_mul3/_073_ ;
 wire \uut.mod_inv.mod_mul3/_074_ ;
 wire \uut.mod_inv.mod_mul3/_075_ ;
 wire \uut.mod_inv.mod_mul3/_076_ ;
 wire \uut.mod_inv.mod_mul3/_077_ ;
 wire \uut.mod_inv.mod_mul3/_078_ ;
 wire \uut.mod_inv.mod_mul3/_079_ ;
 wire \uut.mod_inv.mod_mul3/_080_ ;
 wire \uut.mod_inv.mod_mul3/_081_ ;
 wire \uut.mod_inv.mod_mul3/_082_ ;
 wire \uut.mod_inv.mod_mul3/_083_ ;
 wire \uut.mod_inv.mod_mul3/_084_ ;
 wire \uut.mod_inv.mod_mul3/_085_ ;
 wire \uut.mod_inv.mod_mul3/_086_ ;
 wire \uut.mod_inv.mod_mul3/_087_ ;
 wire \uut.mod_inv.mod_mul3/_088_ ;
 wire \uut.mod_inv.mod_mul3/_089_ ;
 wire \uut.mod_inv.mod_mul3/_090_ ;
 wire \uut.mod_inv.mod_mul3/_091_ ;
 wire \uut.mod_inv.mod_mul3/_092_ ;
 wire \uut.mod_inv.mod_mul3/_093_ ;
 wire \uut.mod_inv.mod_mul3/_094_ ;
 wire \uut.mod_inv.mod_mul3/_095_ ;
 wire \uut.mod_inv.mod_mul3/_096_ ;
 wire \uut.mod_inv.mod_mul3/_097_ ;
 wire \uut.mod_inv.mod_mul3/_098_ ;
 wire \uut.mod_inv.mod_mul3/_099_ ;
 wire \uut.mod_inv.mod_mul3/_100_ ;
 wire \uut.mod_inv.mod_mul3/_101_ ;
 wire \uut.mod_inv.mod_mul3/_102_ ;
 wire \uut.mod_inv.mod_mul3/_103_ ;
 wire \uut.mod_inv.mod_mul3/_104_ ;
 wire \uut.mod_inv.mod_mul3/_105_ ;
 wire \uut.mod_inv.mod_mul3/_106_ ;
 wire \uut.mod_inv.mod_mul3/_107_ ;
 wire \uut.mod_inv.mod_mul3/_108_ ;
 wire \uut.mod_inv.mod_mul3/_109_ ;
 wire \uut.mod_inv.mod_mul3/_110_ ;
 wire \uut.mod_inv.mod_mul3/_111_ ;
 wire \uut.mod_inv.mod_mul3/_112_ ;
 wire \uut.mod_inv.mod_mul3/_113_ ;
 wire \uut.mod_inv.mod_mul3/_114_ ;
 wire \uut.mod_inv.mod_mul3/_115_ ;
 wire \uut.mod_inv.mod_mul3/_116_ ;
 wire \uut.mod_inv.mod_mul3/_117_ ;
 wire \uut.mod_inv.mod_mul3/_118_ ;
 wire \uut.mod_inv.mod_mul3/_119_ ;
 wire \uut.mod_inv.mod_mul3/_120_ ;
 wire \uut.mod_inv.mod_mul3/_121_ ;
 wire \uut.mod_inv.mod_mul3/_122_ ;
 wire \uut.mod_inv.mod_mul3/_123_ ;
 wire \uut.mod_inv.mod_mul3/_124_ ;
 wire \uut.mod_inv.mod_mul3/_125_ ;
 wire \uut.mod_inv.mod_mul3/_126_ ;
 wire \uut.mod_inv.mod_mul3/_127_ ;
 wire \uut.mod_inv.mod_mul3/_128_ ;
 wire \uut.mod_inv.mod_mul3/_129_ ;
 wire \uut.mod_inv.mod_mul3/_130_ ;
 wire \uut.mod_inv.mod_mul3/_131_ ;
 wire \uut.mod_inv.mod_mul3/_132_ ;
 wire \uut.mod_inv.mod_mul3/_133_ ;
 wire \uut.mod_inv.mod_mul3/_134_ ;
 wire \uut.mod_inv.mod_mul3/_135_ ;
 wire \uut.mod_inv.mod_mul3/_136_ ;
 wire \uut.mod_inv.mod_mul3/_137_ ;
 wire \uut.mod_inv.mod_mul3/_138_ ;
 wire \uut.mod_inv.mod_mul3/_139_ ;
 wire \uut.mod_inv.mod_mul3/_140_ ;
 wire \uut.mod_inv.mod_mul3/_141_ ;
 wire \uut.mod_inv.mod_mul3/_142_ ;
 wire \uut.mod_inv.mod_mul3/_143_ ;
 wire \uut.mod_inv.mod_mul3/_144_ ;
 wire \uut.mod_inv.mod_mul3/_145_ ;
 wire \uut.mod_inv.mod_mul3/_146_ ;
 wire \uut.mod_inv.mod_mul3/_147_ ;
 wire \uut.mod_inv.mod_mul3/_148_ ;
 wire \uut.mod_inv.mod_mul3/_149_ ;
 wire \uut.mod_inv.mod_mul3/_150_ ;
 wire \uut.mod_inv.mod_mul3/_151_ ;
 wire \uut.mod_inv.mod_mul3/_152_ ;
 wire \uut.mod_inv.mod_mul3/_153_ ;
 wire \uut.mod_inv.mod_mul3/_154_ ;
 wire \uut.mod_inv.mod_mul3/_155_ ;
 wire \uut.mod_inv.mod_mul3/_156_ ;
 wire \uut.mod_inv.mod_mul3/_157_ ;
 wire \uut.mod_inv.mod_mul3/_158_ ;
 wire \uut.mod_inv.mod_mul3/_159_ ;
 wire \uut.mod_inv.mod_mul3/_160_ ;
 wire \uut.mod_inv.mod_mul3/_161_ ;
 wire \uut.mod_inv.mod_mul3/_162_ ;
 wire \uut.mod_inv.mod_mul3/_163_ ;
 wire \uut.mod_inv.mod_mul3/_164_ ;
 wire \uut.mod_inv.mod_mul3/_165_ ;
 wire \uut.mod_inv.mod_mul3/_166_ ;
 wire \uut.mod_inv.mod_mul3/_167_ ;
 wire \uut.mod_inv.mod_mul3/_168_ ;
 wire \uut.mod_inv.mod_mul3/_169_ ;
 wire \uut.mod_inv.mod_mul3/_170_ ;
 wire \uut.mod_inv.mod_mul3/_171_ ;
 wire \uut.mod_inv.mod_mul3/_172_ ;
 wire \uut.mod_inv.mod_mul3/_173_ ;
 wire \uut.mod_inv.mod_mul3/_174_ ;
 wire \uut.mod_inv.mod_mul3/_175_ ;
 wire \uut.mod_inv.mod_mul3/_176_ ;
 wire \uut.mod_inv.mod_mul3/_177_ ;
 wire \uut.mod_inv.mod_mul3/_178_ ;
 wire \uut.mod_inv.mod_mul3/_179_ ;
 wire \uut.mod_inv.mod_mul3/_180_ ;
 wire \uut.mod_inv.mod_mul3/_181_ ;
 wire \uut.mod_inv.mod_mul3/_182_ ;
 wire \uut.mod_inv.mod_mul3/_183_ ;
 wire \uut.mod_inv.mod_mul3/_184_ ;
 wire \uut.mod_inv.mod_mul3/_185_ ;
 wire \uut.mod_inv.mod_mul3/_186_ ;
 wire \uut.mod_inv.mod_mul3/_187_ ;
 wire \uut.mod_inv.mod_mul3/_188_ ;
 wire \uut.mod_inv.mod_mul3/_189_ ;
 wire \uut.mod_inv.mod_mul3/_190_ ;
 wire \uut.mod_inv.mod_mul3/_191_ ;
 wire \uut.mod_inv.mod_mul3/_192_ ;
 wire \uut.mod_inv.mod_mul3/_193_ ;
 wire \uut.mod_inv.mod_mul3/_194_ ;
 wire \uut.mod_inv.mod_mul3/_195_ ;
 wire \uut.mod_inv.mod_mul3/_196_ ;
 wire \uut.mod_inv.mod_mul3/_197_ ;
 wire \uut.mod_inv.mod_mul3/_198_ ;
 wire \uut.mod_inv.mod_mul3/_199_ ;
 wire \uut.mod_inv.mod_mul3/_200_ ;
 wire \uut.mod_inv.mod_mul3/_201_ ;
 wire \uut.mod_inv.mod_mul3/_202_ ;
 wire \uut.mod_inv.mod_mul3/_203_ ;
 wire \uut.mod_inv.mod_mul3/_204_ ;
 wire \uut.mod_inv.mod_mul3/_205_ ;
 wire \uut.mod_inv.mod_mul3/_206_ ;
 wire \uut.mod_inv.mod_mul3/_207_ ;
 wire \uut.mod_inv.mod_mul3/_208_ ;
 wire \uut.mod_inv.mod_mul3/_209_ ;
 wire \uut.mod_inv.mod_mul3/_210_ ;
 wire \uut.mod_inv.mod_mul3/_211_ ;
 wire \uut.mod_inv.mod_mul3/_212_ ;
 wire \uut.mod_inv.mod_mul3/_213_ ;
 wire \uut.mod_inv.mod_mul3/_214_ ;
 wire \uut.mod_inv.mod_mul3/_215_ ;
 wire \uut.mod_inv.mod_mul3/_216_ ;
 wire \uut.mod_inv.mod_mul3/_217_ ;
 wire \uut.mod_inv.mod_mul3/_218_ ;
 wire \uut.mod_inv.mod_mul3/_219_ ;
 wire \uut.mod_inv.mod_mul3/_220_ ;
 wire \uut.mod_inv.mod_mul3_out1[0] ;
 wire \uut.mod_inv.mod_mul3_out1[1] ;
 wire \uut.mod_inv.mod_mul3_out1[2] ;
 wire \uut.mod_inv.mod_mul3_out1[3] ;
 wire \uut.mod_inv.mod_mul3_out2[0] ;
 wire \uut.mod_inv.mod_mul3_out2[1] ;
 wire \uut.mod_inv.mod_mul3_out2[2] ;
 wire \uut.mod_inv.mod_mul3_out2[3] ;
 wire \uut.mod_inv.mod_mul3_out3[0] ;
 wire \uut.mod_inv.mod_mul3_out3[1] ;
 wire \uut.mod_inv.mod_mul3_out3[2] ;
 wire \uut.mod_inv.mod_mul3_out3[3] ;
 wire \uut.mod_inv.mul_in1[0] ;
 wire \uut.mod_inv.mul_in1[1] ;
 wire \uut.mod_inv.mul_in1[2] ;
 wire \uut.mod_inv.mul_in1[3] ;
 wire \uut.mod_inv.mul_in3[0] ;
 wire \uut.mod_inv.mul_in3[1] ;
 wire \uut.mod_inv.mul_in3[2] ;
 wire \uut.mod_inv.mul_in3[3] ;
 wire \uut.mod_inv.random_xor_1[0] ;
 wire \uut.mod_inv.random_xor_1[1] ;
 wire \uut.mod_inv.random_xor_1[2] ;
 wire \uut.mod_inv.random_xor_1[3] ;
 wire \uut.mod_inv.random_xor_2[0] ;
 wire \uut.mod_inv.random_xor_2[1] ;
 wire \uut.mod_inv.random_xor_2[2] ;
 wire \uut.mod_inv.random_xor_2[3] ;
 wire \uut.mod_inv.sh1_reg_0_1[0] ;
 wire \uut.mod_inv.sh1_reg_0_1[1] ;
 wire \uut.mod_inv.sh1_reg_0_1[2] ;
 wire \uut.mod_inv.sh1_reg_0_1[3] ;
 wire \uut.mod_inv.sh1_reg_0_2[0] ;
 wire \uut.mod_inv.sh1_reg_0_2[1] ;
 wire \uut.mod_inv.sh1_reg_0_2[2] ;
 wire \uut.mod_inv.sh1_reg_0_2[3] ;
 wire \uut.mod_inv.sh1_reg_1_1[0] ;
 wire \uut.mod_inv.sh1_reg_1_1[1] ;
 wire \uut.mod_inv.sh1_reg_1_1[2] ;
 wire \uut.mod_inv.sh1_reg_1_1[3] ;
 wire \uut.mod_inv.sh1_reg_1_2[0] ;
 wire \uut.mod_inv.sh1_reg_1_2[1] ;
 wire \uut.mod_inv.sh1_reg_1_2[2] ;
 wire \uut.mod_inv.sh1_reg_1_2[3] ;
 wire \uut.mod_inv.sh1_xor_out[0] ;
 wire \uut.mod_inv.sh1_xor_out[1] ;
 wire \uut.mod_inv.sh1_xor_out[2] ;
 wire \uut.mod_inv.sh1_xor_out[3] ;
 wire \uut.mod_inv.sh2_reg_0_1[0] ;
 wire \uut.mod_inv.sh2_reg_0_1[1] ;
 wire \uut.mod_inv.sh2_reg_0_1[2] ;
 wire \uut.mod_inv.sh2_reg_0_1[3] ;
 wire \uut.mod_inv.sh2_reg_0_2[0] ;
 wire \uut.mod_inv.sh2_reg_0_2[1] ;
 wire \uut.mod_inv.sh2_reg_0_2[2] ;
 wire \uut.mod_inv.sh2_reg_0_2[3] ;
 wire \uut.mod_inv.sh2_reg_1_1[0] ;
 wire \uut.mod_inv.sh2_reg_1_1[1] ;
 wire \uut.mod_inv.sh2_reg_1_1[2] ;
 wire \uut.mod_inv.sh2_reg_1_1[3] ;
 wire \uut.mod_inv.sh2_reg_1_2[0] ;
 wire \uut.mod_inv.sh2_reg_1_2[1] ;
 wire \uut.mod_inv.sh2_reg_1_2[2] ;
 wire \uut.mod_inv.sh2_reg_1_2[3] ;
 wire \uut.mod_inv.sh3_reg_0_1[0] ;
 wire \uut.mod_inv.sh3_reg_0_1[1] ;
 wire \uut.mod_inv.sh3_reg_0_1[2] ;
 wire \uut.mod_inv.sh3_reg_0_1[3] ;
 wire \uut.mod_inv.sh3_reg_0_2[0] ;
 wire \uut.mod_inv.sh3_reg_0_2[1] ;
 wire \uut.mod_inv.sh3_reg_0_2[2] ;
 wire \uut.mod_inv.sh3_reg_0_2[3] ;
 wire \uut.mod_inv.sh3_reg_1_1[0] ;
 wire \uut.mod_inv.sh3_reg_1_1[1] ;
 wire \uut.mod_inv.sh3_reg_1_1[2] ;
 wire \uut.mod_inv.sh3_reg_1_1[3] ;
 wire \uut.mod_inv.sh3_reg_1_2[0] ;
 wire \uut.mod_inv.sh3_reg_1_2[1] ;
 wire \uut.mod_inv.sh3_reg_1_2[2] ;
 wire \uut.mod_inv.sh3_reg_1_2[3] ;
 wire \uut.mod_inv.sq_scl_in[0] ;
 wire \uut.mod_inv.sq_scl_in[1] ;
 wire \uut.mod_inv.sq_scl_in[2] ;
 wire \uut.mod_inv.sq_scl_in[3] ;
 wire \uut.mod_inv.sq_scl_out1[0] ;
 wire \uut.mod_inv.sq_scl_out1[1] ;
 wire \uut.mod_inv.sq_scl_out1[2] ;
 wire \uut.mod_inv.sq_scl_out1[3] ;
 wire \uut.mod_inv.sq_scl_out2[0] ;
 wire \uut.mod_inv.sq_scl_out2[1] ;
 wire \uut.mod_inv.sq_scl_out2[2] ;
 wire \uut.mod_inv.sq_scl_out2[3] ;
 wire \uut.mod_inv.sq_scl_out2_reg[0] ;
 wire \uut.mod_inv.sq_scl_out2_reg[1] ;
 wire \uut.mod_inv.sq_scl_out2_reg[2] ;
 wire \uut.mod_inv.sq_scl_out2_reg[3] ;
 wire \uut.sel_in_sh1.m0.Q ;
 wire \uut.sel_in_sh1.m1.Q ;
 wire \uut.sel_in_sh1.m3.Q ;
 wire \uut.sel_in_sh1.m4.Q ;
 wire \uut.sel_in_sh1.m5.Q ;
 wire \uut.sel_in_sh1.m6.Q ;
 wire \uut.sel_in_sh1.m7.Q ;
 wire \uut.sel_in_sh2.m0.Q ;
 wire \uut.sel_in_sh2.m1.Q ;
 wire \uut.sel_in_sh2.m3.Q ;
 wire \uut.sel_in_sh2.m4.Q ;
 wire \uut.sel_in_sh2.m5.Q ;
 wire \uut.sel_in_sh2.m6.Q ;
 wire \uut.sel_in_sh2.m7.Q ;
 wire \uut.sel_in_sh3.m0.Q ;
 wire \uut.sel_in_sh3.m1.Q ;
 wire \uut.sel_in_sh3.m3.Q ;
 wire \uut.sel_in_sh3.m4.Q ;
 wire \uut.sel_in_sh3.m5.Q ;
 wire \uut.sel_in_sh3.m6.Q ;
 wire \uut.sel_in_sh3.m7.Q ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\uut.R1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\uut.mod_inv.mul_in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\uut.mod_inv.inv_mod/_244_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_178 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_286 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_180 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_192 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_212 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_228 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_320 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_203 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_215 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_240 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_279 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_330 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_80 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_226 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_288 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_320 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_332 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_182 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_194 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_206 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_214 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_327 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_339 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_328 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_184 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_196 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_208 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_185 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_203 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_265 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_292 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_332 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_200 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_212 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_266 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_204 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_227 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_239 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_336 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_118 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_146 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_232 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_244 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_88 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_182 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_283 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_211 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_256 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_288 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_192 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_204 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_319 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_76 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_124 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_144 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_156 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_282 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_294 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_173 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_238 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_267 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_106 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_170 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_182 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_239 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_94 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_147 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_90 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_128 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_276 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_42 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_34 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_282 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_314 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_326 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_338 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_203 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_260 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_95 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_132 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_260 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_307 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_319 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_184 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_285 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_323 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_335 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_288 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_300 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_312 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_163 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_268 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_50 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_136 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_154 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_77 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_89 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_272 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_338 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_184 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_266 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_297 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_319 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_71 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_103 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_115 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_127 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_45 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_118 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_24 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_98 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_13 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_62 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_140 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_152 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_196 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_255 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_267 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_161 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_228 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_274 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_286 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_263 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_339 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_16 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_202 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_312 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_324 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_71 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_203 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_230 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_191 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_75 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_112 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_146 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_167 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_179 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_215 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_239 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_260 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_272 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_284 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_296 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_318 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_56 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_68 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_116 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_151 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_28 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_10 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_117 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_338 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_129 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_257 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_80 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_184 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_239 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_326 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_338 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_143 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_16 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_209 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_243 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_259 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_28 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_40 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_76 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_203 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_110 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_122 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_16 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_166 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_276 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_288 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_122 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_134 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_146 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_176 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_99 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_326 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_338 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_96 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_214 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_51 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_257 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_107 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_278 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_290 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_328 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_63 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_152 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_191 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_25 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_110 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_122 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_154 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_331 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_237 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_269 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_291 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_40 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_250 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_43 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_100 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_213 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_66 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_88 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_18 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_285 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_297 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_114 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_126 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_323 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_335 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_72 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_244 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_256 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_26 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_323 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_38 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_160 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_62 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_179 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_119 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_286 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_296 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_308 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_320 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_43 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_90 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_189 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_201 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_302 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_314 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_152 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_229 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_323 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_271 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_242 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_254 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_266 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__xor2_4 _0433_ (.A(\uut.in3[6] ),
    .B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__xnor2_4 _0434_ (.A(\uut.in3[1] ),
    .B(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0146_));
 sky130_fd_sc_hd__xor2_4 _0435_ (.A(\uut.in3[7] ),
    .B(\uut.in3[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__xor2_2 _0436_ (.A(\uut.in3[2] ),
    .B(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__xnor2_4 _0437_ (.A(_0146_),
    .B(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh3.m7.Q ));
 sky130_fd_sc_hd__xnor2_4 _0438_ (.A(\uut.in3[5] ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0149_));
 sky130_fd_sc_hd__clkinv_4 _0439_ (.A(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh3.m1.Q ));
 sky130_fd_sc_hd__xnor2_4 _0440_ (.A(\uut.in3[4] ),
    .B(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh3.m6.Q ));
 sky130_fd_sc_hd__xnor2_4 _0441_ (.A(\uut.in3[1] ),
    .B(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh3.m5.Q ));
 sky130_fd_sc_hd__xor2_4 _0442_ (.A(net21),
    .B(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.sel_in_sh3.m4.Q ));
 sky130_fd_sc_hd__xor2_2 _0443_ (.A(\uut.in3[4] ),
    .B(\uut.in3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__xor2_1 _0444_ (.A(\uut.in3[7] ),
    .B(\uut.in3[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__xnor2_2 _0445_ (.A(\uut.in3[0] ),
    .B(_0151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0152_));
 sky130_fd_sc_hd__xnor2_4 _0446_ (.A(_0150_),
    .B(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh3.m3.Q ));
 sky130_fd_sc_hd__xor2_2 _0447_ (.A(\uut.in3[3] ),
    .B(\uut.in3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__xnor2_4 _0448_ (.A(_0146_),
    .B(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh3.m0.Q ));
 sky130_fd_sc_hd__xor2_4 _0449_ (.A(\uut.in2[6] ),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__xnor2_4 _0450_ (.A(\uut.in2[5] ),
    .B(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0155_));
 sky130_fd_sc_hd__xnor2_2 _0451_ (.A(\uut.in2[7] ),
    .B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m4.Q ));
 sky130_fd_sc_hd__xnor2_2 _0452_ (.A(\uut.in2[2] ),
    .B(\uut.in2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0156_));
 sky130_fd_sc_hd__xnor2_4 _0453_ (.A(net12),
    .B(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m7.Q ));
 sky130_fd_sc_hd__inv_2 _0454_ (.A(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m1.Q ));
 sky130_fd_sc_hd__xnor2_4 _0455_ (.A(\uut.in2[4] ),
    .B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m6.Q ));
 sky130_fd_sc_hd__xnor2_4 _0456_ (.A(\uut.in2[1] ),
    .B(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m5.Q ));
 sky130_fd_sc_hd__xnor2_4 _0457_ (.A(\uut.in2[3] ),
    .B(\uut.in2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0157_));
 sky130_fd_sc_hd__xnor2_1 _0458_ (.A(\uut.in2[4] ),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0158_));
 sky130_fd_sc_hd__xnor2_2 _0459_ (.A(\uut.in2[7] ),
    .B(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0159_));
 sky130_fd_sc_hd__xnor2_4 _0460_ (.A(_0157_),
    .B(_0159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m3.Q ));
 sky130_fd_sc_hd__xor2_2 _0461_ (.A(\uut.in2[2] ),
    .B(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__xnor2_4 _0462_ (.A(_0157_),
    .B(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh2.m0.Q ));
 sky130_fd_sc_hd__xor2_4 _0463_ (.A(\uut.in1[6] ),
    .B(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__xnor2_4 _0464_ (.A(\uut.in1[5] ),
    .B(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0162_));
 sky130_fd_sc_hd__xnor2_4 _0465_ (.A(\uut.in1[7] ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m4.Q ));
 sky130_fd_sc_hd__xnor2_2 _0466_ (.A(\uut.in1[2] ),
    .B(\uut.in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0163_));
 sky130_fd_sc_hd__xnor2_4 _0467_ (.A(net11),
    .B(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m7.Q ));
 sky130_fd_sc_hd__inv_2 _0468_ (.A(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m1.Q ));
 sky130_fd_sc_hd__xnor2_4 _0469_ (.A(\uut.in1[4] ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m6.Q ));
 sky130_fd_sc_hd__xnor2_4 _0470_ (.A(\uut.in1[1] ),
    .B(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m5.Q ));
 sky130_fd_sc_hd__xor2_4 _0471_ (.A(\uut.in1[3] ),
    .B(\uut.in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__xor2_2 _0472_ (.A(\uut.in1[4] ),
    .B(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__xnor2_2 _0473_ (.A(\uut.in1[7] ),
    .B(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0166_));
 sky130_fd_sc_hd__xnor2_4 _0474_ (.A(_0164_),
    .B(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m3.Q ));
 sky130_fd_sc_hd__xnor2_2 _0475_ (.A(\uut.in1[2] ),
    .B(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0167_));
 sky130_fd_sc_hd__xnor2_4 _0476_ (.A(_0164_),
    .B(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.sel_in_sh1.m0.Q ));
 sky130_fd_sc_hd__xor2_2 _0477_ (.A(\uut.sel_in_sh1.m4.Q ),
    .B(\uut.sel_in_sh1.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sh1_xor_out[0] ));
 sky130_fd_sc_hd__clkbuf_1 _0478_ (.A(\uut.in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__buf_1 _0479_ (.A(_0168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sh1_xor_out[1] ));
 sky130_fd_sc_hd__xnor2_1 _0480_ (.A(net95),
    .B(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.sh1_xor_out[2] ));
 sky130_fd_sc_hd__xor2_1 _0481_ (.A(\uut.sel_in_sh1.m7.Q ),
    .B(\uut.sel_in_sh1.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sh1_xor_out[3] ));
 sky130_fd_sc_hd__xnor2_1 _0482_ (.A(\uut.sel_in_sh3.m4.Q ),
    .B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0169_));
 sky130_fd_sc_hd__xor2_1 _0483_ (.A(\uut.sel_in_sh3.m0.Q ),
    .B(\uut.sel_in_sh2.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__xnor2_2 _0484_ (.A(_0169_),
    .B(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.sq_scl_in[0] ));
 sky130_fd_sc_hd__xor2_2 _0485_ (.A(\uut.in2[1] ),
    .B(\uut.in3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_in[1] ));
 sky130_fd_sc_hd__xor2_1 _0486_ (.A(net27),
    .B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__xnor2_1 _0487_ (.A(\uut.sel_in_sh3.m6.Q ),
    .B(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0172_));
 sky130_fd_sc_hd__xnor2_1 _0488_ (.A(\uut.sel_in_sh2.m6.Q ),
    .B(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.sq_scl_in[2] ));
 sky130_fd_sc_hd__xor2_1 _0489_ (.A(\uut.sel_in_sh3.m7.Q ),
    .B(\uut.sel_in_sh3.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__xnor2_1 _0490_ (.A(\uut.sel_in_sh2.m7.Q ),
    .B(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0174_));
 sky130_fd_sc_hd__xnor2_1 _0491_ (.A(\uut.sel_in_sh2.m3.Q ),
    .B(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.sq_scl_in[3] ));
 sky130_fd_sc_hd__xor2_4 _0492_ (.A(\uut.mod_inv.random_xor_1[0] ),
    .B(\uut.mod_inv.sq_scl_out2_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in2[0] ));
 sky130_fd_sc_hd__xor2_2 _0493_ (.A(\uut.mod_inv.random_xor_1[1] ),
    .B(\uut.mod_inv.sq_scl_out2_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in2[1] ));
 sky130_fd_sc_hd__xor2_4 _0494_ (.A(\uut.mod_inv.random_xor_1[2] ),
    .B(\uut.mod_inv.sq_scl_out2_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in2[2] ));
 sky130_fd_sc_hd__xor2_2 _0495_ (.A(\uut.mod_inv.random_xor_1[3] ),
    .B(\uut.mod_inv.sq_scl_out2_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in2[3] ));
 sky130_fd_sc_hd__xor2_4 _0496_ (.A(\uut.mod_inv.mod_mul1_out2_xor[0] ),
    .B(\uut.mod_inv.mod_mul1_out1_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in3[0] ));
 sky130_fd_sc_hd__xor2_4 _0497_ (.A(\uut.mod_inv.mod_mul1_out2_xor[1] ),
    .B(\uut.mod_inv.mod_mul1_out1_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in3[1] ));
 sky130_fd_sc_hd__xor2_1 _0498_ (.A(\uut.mod_inv.mod_mul1_out2_xor[2] ),
    .B(\uut.mod_inv.mod_mul1_out1_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in3[2] ));
 sky130_fd_sc_hd__xor2_4 _0499_ (.A(\uut.mod_inv.mod_mul1_out2_xor[3] ),
    .B(\uut.mod_inv.mod_mul1_out1_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_in3[3] ));
 sky130_fd_sc_hd__xor2_4 _0500_ (.A(\uut.mod_inv.inv_out2_xor[0] ),
    .B(\uut.mod_inv.inv_out1_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in1[0] ));
 sky130_fd_sc_hd__xor2_2 _0501_ (.A(\uut.mod_inv.inv_out2_xor[1] ),
    .B(\uut.mod_inv.inv_out1_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in1[1] ));
 sky130_fd_sc_hd__xor2_4 _0502_ (.A(\uut.mod_inv.inv_out2_xor[2] ),
    .B(\uut.mod_inv.inv_out1_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in1[2] ));
 sky130_fd_sc_hd__xor2_4 _0503_ (.A(\uut.mod_inv.inv_out2_xor[3] ),
    .B(\uut.mod_inv.inv_out1_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in1[3] ));
 sky130_fd_sc_hd__xor2_2 _0504_ (.A(\uut.mod_inv.random_xor_2[0] ),
    .B(\uut.mod_inv.inv_out4_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in3[0] ));
 sky130_fd_sc_hd__xor2_2 _0505_ (.A(\uut.mod_inv.random_xor_2[1] ),
    .B(\uut.mod_inv.inv_out4_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in3[1] ));
 sky130_fd_sc_hd__xor2_2 _0506_ (.A(\uut.mod_inv.random_xor_2[2] ),
    .B(\uut.mod_inv.inv_out4_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in3[2] ));
 sky130_fd_sc_hd__xor2_4 _0507_ (.A(\uut.mod_inv.random_xor_2[3] ),
    .B(\uut.mod_inv.inv_out4_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mul_in3[3] ));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0175_));
 sky130_fd_sc_hd__buf_4 _0509_ (.A(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__a21oi_1 _0510_ (.A1(\uut.R0[4] ),
    .A2(\uut.R0[0] ),
    .B1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0177_));
 sky130_fd_sc_hd__o21a_1 _0511_ (.A1(\uut.R0[4] ),
    .A2(net72),
    .B1(_0177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0000_));
 sky130_fd_sc_hd__a21oi_1 _0512_ (.A1(\uut.R0[5] ),
    .A2(\uut.R0[1] ),
    .B1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0178_));
 sky130_fd_sc_hd__o21a_1 _0513_ (.A1(\uut.R0[5] ),
    .A2(net76),
    .B1(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__a21oi_1 _0514_ (.A1(\uut.R0[6] ),
    .A2(\uut.R0[2] ),
    .B1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0179_));
 sky130_fd_sc_hd__o21a_1 _0515_ (.A1(\uut.R0[6] ),
    .A2(net85),
    .B1(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _0516_ (.A(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__a21oi_1 _0517_ (.A1(\uut.R0[7] ),
    .A2(\uut.R0[3] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0181_));
 sky130_fd_sc_hd__o21a_1 _0518_ (.A1(\uut.R0[7] ),
    .A2(net74),
    .B1(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0003_));
 sky130_fd_sc_hd__buf_2 _0519_ (.A(\out_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__or2_2 _0520_ (.A(\out_count[1] ),
    .B(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__xor2_2 _0521_ (.A(\uut.mod_inv.mod_mul3_out2[2] ),
    .B(\uut.mod_inv.mod_mul3_out2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__or2_1 _0522_ (.A(\uut.mod_inv.mod_mul2_out2[1] ),
    .B(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__nand2_1 _0523_ (.A(\uut.mod_inv.mod_mul2_out2[1] ),
    .B(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0186_));
 sky130_fd_sc_hd__a31o_1 _0524_ (.A1(\out_count[1] ),
    .A2(_0185_),
    .A3(_0186_),
    .B1(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_1 _0525_ (.A(\out_count[1] ),
    .B(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0188_));
 sky130_fd_sc_hd__xnor2_2 _0526_ (.A(\uut.mod_inv.mod_mul3_out3[2] ),
    .B(\uut.mod_inv.mod_mul3_out3[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0189_));
 sky130_fd_sc_hd__xnor2_1 _0527_ (.A(\uut.mod_inv.mod_mul2_out3[1] ),
    .B(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0190_));
 sky130_fd_sc_hd__xnor2_1 _0528_ (.A(\uut.mod_inv.mod_mul3_out1[2] ),
    .B(\uut.mod_inv.mod_mul3_out1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0191_));
 sky130_fd_sc_hd__xnor2_1 _0529_ (.A(\uut.mod_inv.mod_mul2_out1[1] ),
    .B(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0192_));
 sky130_fd_sc_hd__o22a_1 _0530_ (.A1(_0188_),
    .A2(_0190_),
    .B1(_0192_),
    .B2(\out_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__nand2_1 _0531_ (.A(_0187_),
    .B(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0194_));
 sky130_fd_sc_hd__clkbuf_4 _0532_ (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _0533_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__o211a_1 _0534_ (.A1(uo_out[0]),
    .A2(_0183_),
    .B1(_0194_),
    .C1(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(\out_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0197_));
 sky130_fd_sc_hd__nand2_1 _0536_ (.A(_0197_),
    .B(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0198_));
 sky130_fd_sc_hd__xor2_1 _0537_ (.A(\uut.mod_inv.mod_mul2_out1[1] ),
    .B(\uut.mod_inv.mod_mul3_out1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_1 _0538_ (.A(\uut.mod_inv.mod_mul3_out1[0] ),
    .B(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0200_));
 sky130_fd_sc_hd__xor2_1 _0539_ (.A(\uut.mod_inv.mod_mul2_out3[1] ),
    .B(\uut.mod_inv.mod_mul3_out3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__xnor2_1 _0540_ (.A(\uut.mod_inv.mod_mul3_out3[0] ),
    .B(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0202_));
 sky130_fd_sc_hd__clkbuf_4 _0541_ (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__o221a_1 _0542_ (.A1(uo_out[1]),
    .A2(_0183_),
    .B1(_0202_),
    .B2(_0188_),
    .C1(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__xnor2_1 _0543_ (.A(\uut.mod_inv.mod_mul3_out2[0] ),
    .B(\uut.mod_inv.mod_mul2_out2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0205_));
 sky130_fd_sc_hd__or2_1 _0544_ (.A(\uut.mod_inv.mod_mul3_out2[1] ),
    .B(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _0545_ (.A(\uut.mod_inv.mod_mul3_out2[1] ),
    .B(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0207_));
 sky130_fd_sc_hd__or2_2 _0546_ (.A(_0197_),
    .B(\out_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__a21o_1 _0547_ (.A1(_0206_),
    .A2(_0207_),
    .B1(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0209_));
 sky130_fd_sc_hd__o211a_1 _0548_ (.A1(_0198_),
    .A2(_0200_),
    .B1(_0204_),
    .C1(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0005_));
 sky130_fd_sc_hd__xnor2_2 _0549_ (.A(\uut.mod_inv.mod_mul3_out3[1] ),
    .B(\uut.mod_inv.mod_mul2_out3[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0210_));
 sky130_fd_sc_hd__xor2_1 _0550_ (.A(\uut.mod_inv.mod_mul3_out3[2] ),
    .B(\uut.mod_inv.mod_mul2_out3[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__xnor2_1 _0551_ (.A(\uut.mod_inv.mod_mul2_out3[2] ),
    .B(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0212_));
 sky130_fd_sc_hd__xnor2_1 _0552_ (.A(_0210_),
    .B(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0213_));
 sky130_fd_sc_hd__xor2_2 _0553_ (.A(\uut.mod_inv.mod_mul3_out2[1] ),
    .B(\uut.mod_inv.mod_mul2_out2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__xor2_1 _0554_ (.A(\uut.mod_inv.mod_mul3_out2[2] ),
    .B(\uut.mod_inv.mod_mul2_out2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__xnor2_1 _0555_ (.A(\uut.mod_inv.mod_mul2_out2[2] ),
    .B(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0216_));
 sky130_fd_sc_hd__a21o_1 _0556_ (.A1(_0214_),
    .A2(_0216_),
    .B1(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__nor2_1 _0557_ (.A(_0214_),
    .B(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0218_));
 sky130_fd_sc_hd__o2bb2a_1 _0558_ (.A1_N(_0208_),
    .A2_N(_0213_),
    .B1(_0217_),
    .B2(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__xor2_2 _0559_ (.A(\uut.mod_inv.mod_mul3_out1[2] ),
    .B(\uut.mod_inv.mod_mul2_out1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__xnor2_2 _0560_ (.A(\uut.mod_inv.mod_mul3_out1[1] ),
    .B(\uut.mod_inv.mod_mul2_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0221_));
 sky130_fd_sc_hd__xor2_1 _0561_ (.A(\uut.mod_inv.mod_mul2_out1[2] ),
    .B(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__nor2_1 _0562_ (.A(_0220_),
    .B(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0223_));
 sky130_fd_sc_hd__a21o_1 _0563_ (.A1(_0220_),
    .A2(_0222_),
    .B1(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__o221a_1 _0564_ (.A1(uo_out[2]),
    .A2(_0183_),
    .B1(_0223_),
    .B2(_0224_),
    .C1(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__o21a_1 _0565_ (.A1(_0197_),
    .A2(_0219_),
    .B1(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0006_));
 sky130_fd_sc_hd__xnor2_1 _0566_ (.A(\uut.mod_inv.mod_mul3_out2[3] ),
    .B(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _0567_ (.A(_0184_),
    .B(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ba_1 _0568_ (.A1(_0184_),
    .A2(_0226_),
    .B1_N(\out_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__xnor2_1 _0569_ (.A(\uut.mod_inv.mod_mul3_out3[3] ),
    .B(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0229_));
 sky130_fd_sc_hd__xor2_1 _0570_ (.A(_0189_),
    .B(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__a221o_1 _0571_ (.A1(_0227_),
    .A2(_0228_),
    .B1(_0230_),
    .B2(_0182_),
    .C1(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _0572_ (.A(\out_count[1] ),
    .B(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _0573_ (.A(net94),
    .B(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0233_));
 sky130_fd_sc_hd__xnor2_1 _0574_ (.A(\uut.mod_inv.mod_mul3_out1[3] ),
    .B(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _0575_ (.A(_0191_),
    .B(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0235_));
 sky130_fd_sc_hd__or2_1 _0576_ (.A(_0191_),
    .B(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__a21o_1 _0577_ (.A1(_0235_),
    .A2(_0236_),
    .B1(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__a31oi_1 _0578_ (.A1(_0231_),
    .A2(_0233_),
    .A3(_0237_),
    .B1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0007_));
 sky130_fd_sc_hd__and2_1 _0579_ (.A(_0197_),
    .B(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _0580_ (.A1(uo_out[4]),
    .A2(_0232_),
    .B1(_0238_),
    .B2(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__and3_1 _0581_ (.A(\out_count[1] ),
    .B(_0182_),
    .C(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_1 _0582_ (.A(_0208_),
    .B(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0241_));
 sky130_fd_sc_hd__o31a_1 _0583_ (.A1(_0239_),
    .A2(_0240_),
    .A3(_0241_),
    .B1(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__o2bb2a_1 _0584_ (.A1_N(uo_out[5]),
    .A2_N(_0232_),
    .B1(_0198_),
    .B2(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__o22a_1 _0585_ (.A1(_0208_),
    .A2(_0215_),
    .B1(_0211_),
    .B2(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__a21oi_1 _0586_ (.A1(_0242_),
    .A2(_0243_),
    .B1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0009_));
 sky130_fd_sc_hd__xnor2_1 _0587_ (.A(\uut.mod_inv.mod_mul2_out2[3] ),
    .B(\uut.mod_inv.mod_mul3_out2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0244_));
 sky130_fd_sc_hd__xnor2_1 _0588_ (.A(\uut.mod_inv.mod_mul2_out1[3] ),
    .B(\uut.mod_inv.mod_mul3_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0245_));
 sky130_fd_sc_hd__xnor2_1 _0589_ (.A(\uut.mod_inv.mod_mul2_out3[3] ),
    .B(\uut.mod_inv.mod_mul3_out3[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0246_));
 sky130_fd_sc_hd__mux4_1 _0590_ (.A0(uo_out[6]),
    .A1(_0244_),
    .A2(_0245_),
    .A3(_0246_),
    .S0(\out_count[1] ),
    .S1(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__and2_1 _0591_ (.A(_0196_),
    .B(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_1 _0592_ (.A(_0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__a2bb2o_1 _0593_ (.A1_N(_0198_),
    .A2_N(_0221_),
    .B1(uo_out[7]),
    .B2(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_1 _0594_ (.A(_0188_),
    .B(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0250_));
 sky130_fd_sc_hd__and2b_1 _0595_ (.A_N(_0208_),
    .B(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__o31a_1 _0596_ (.A1(_0249_),
    .A2(_0250_),
    .A3(_0251_),
    .B1(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0011_));
 sky130_fd_sc_hd__nand2_1 _0597_ (.A(net83),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0252_));
 sky130_fd_sc_hd__o211a_1 _0598_ (.A1(net83),
    .A2(_0182_),
    .B1(_0196_),
    .C1(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__o211a_1 _0599_ (.A1(net83),
    .A2(net89),
    .B1(_0196_),
    .C1(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _0600_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(\uut.R1[0] ),
    .A1(net3),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__and2_1 _0602_ (.A(_0196_),
    .B(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_1 _0603_ (.A(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(\uut.R1[1] ),
    .A1(net4),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__and2_1 _0605_ (.A(_0196_),
    .B(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_1 _0606_ (.A(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0607_ (.A0(\uut.R1[2] ),
    .A1(net5),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__and2_1 _0608_ (.A(_0196_),
    .B(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _0609_ (.A(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(\uut.R1[3] ),
    .A1(net6),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__and2_1 _0611_ (.A(_0196_),
    .B(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _0613_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(\uut.R1[4] ),
    .A1(net7),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__and2_1 _0615_ (.A(_0262_),
    .B(_0263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0617_ (.A0(\uut.R1[5] ),
    .A1(net8),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__and2_1 _0618_ (.A(_0262_),
    .B(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__clkbuf_1 _0619_ (.A(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0620_ (.A0(\uut.R1[6] ),
    .A1(net9),
    .S(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__and2_1 _0621_ (.A(_0262_),
    .B(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _0622_ (.A(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_4 _0623_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(\uut.R1[7] ),
    .A1(net10),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(_0262_),
    .B(_0270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _0626_ (.A(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(\uut.R0[0] ),
    .A1(\uut.R1[0] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _0628_ (.A(_0262_),
    .B(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _0629_ (.A(_0273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(\uut.R0[1] ),
    .A1(\uut.R1[1] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__and2_1 _0631_ (.A(_0262_),
    .B(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(\uut.R0[2] ),
    .A1(\uut.R1[2] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _0634_ (.A(_0262_),
    .B(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_1 _0635_ (.A(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(\uut.R0[3] ),
    .A1(\uut.R1[3] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__and2_1 _0637_ (.A(_0262_),
    .B(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_1 _0638_ (.A(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(\uut.R0[4] ),
    .A1(\uut.R1[4] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__and2_1 _0640_ (.A(_0262_),
    .B(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _0641_ (.A(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(\uut.R0[5] ),
    .A1(\uut.R1[5] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _0643_ (.A(_0262_),
    .B(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_2 _0645_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(\uut.R0[6] ),
    .A1(\uut.R1[6] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__and2_1 _0647_ (.A(_0284_),
    .B(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(\uut.R0[7] ),
    .A1(\uut.R1[7] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__and2_1 _0650_ (.A(_0284_),
    .B(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(\uut.in3[0] ),
    .A1(\uut.R0[0] ),
    .S(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__and2_1 _0653_ (.A(_0284_),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _0654_ (.A(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_4 _0655_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _0656_ (.A0(\uut.in3[1] ),
    .A1(\uut.R0[1] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__and2_1 _0657_ (.A(_0284_),
    .B(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0658_ (.A(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(\uut.in3[2] ),
    .A1(\uut.R0[2] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__and2_1 _0660_ (.A(_0284_),
    .B(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0661_ (.A(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(\uut.in3[3] ),
    .A1(\uut.R0[3] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__and2_1 _0663_ (.A(_0284_),
    .B(_0296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0665_ (.A0(\uut.in3[4] ),
    .A1(\uut.R0[4] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__and2_1 _0666_ (.A(_0284_),
    .B(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0667_ (.A(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0668_ (.A0(\uut.in3[5] ),
    .A1(\uut.R0[5] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _0669_ (.A(_0284_),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0670_ (.A(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0671_ (.A0(\uut.in3[6] ),
    .A1(\uut.R0[6] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__and2_1 _0672_ (.A(_0284_),
    .B(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _0673_ (.A(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0674_ (.A0(\uut.in3[7] ),
    .A1(\uut.R0[7] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__and2_1 _0675_ (.A(_0284_),
    .B(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _0676_ (.A(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _0677_ (.A(\uut.in3[0] ),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(_0253_),
    .B(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0307_));
 sky130_fd_sc_hd__o22a_1 _0680_ (.A1(_0253_),
    .A2(net92),
    .B1(_0123_),
    .B2(_0307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__buf_2 _0681_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _0682_ (.A0(\uut.in2[1] ),
    .A1(\uut.in3[1] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__and2_1 _0683_ (.A(_0308_),
    .B(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0684_ (.A(_0310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0685_ (.A0(\uut.in2[2] ),
    .A1(\uut.in3[2] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _0686_ (.A(_0308_),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0687_ (.A(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(\uut.in2[3] ),
    .A1(\uut.in3[3] ),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__and2_1 _0689_ (.A(_0308_),
    .B(_0313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0690_ (.A(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__clkbuf_4 _0691_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(\uut.in2[4] ),
    .A1(\uut.in3[4] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__and2_1 _0693_ (.A(_0308_),
    .B(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _0694_ (.A(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(\uut.in2[5] ),
    .A1(\uut.in3[5] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__and2_1 _0696_ (.A(_0308_),
    .B(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(\uut.in2[6] ),
    .A1(\uut.in3[6] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__and2_1 _0699_ (.A(_0308_),
    .B(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0701_ (.A0(\uut.in2[7] ),
    .A1(\uut.in3[7] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _0702_ (.A(_0308_),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _0704_ (.A(\uut.in2[0] ),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _0705_ (.A(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0119_));
 sky130_fd_sc_hd__o22a_1 _0706_ (.A1(_0253_),
    .A2(\uut.in1[0] ),
    .B1(_0307_),
    .B2(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(\uut.in1[1] ),
    .A1(\uut.in2[1] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(_0308_),
    .B(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(\uut.in1[2] ),
    .A1(\uut.in2[2] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(_0308_),
    .B(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(\uut.in1[3] ),
    .A1(\uut.in2[3] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _0714_ (.A(_0308_),
    .B(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0715_ (.A(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__clkbuf_2 _0716_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(\uut.in1[4] ),
    .A1(\uut.in2[4] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _0718_ (.A(_0331_),
    .B(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _0719_ (.A(_0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(\uut.in1[5] ),
    .A1(\uut.in2[5] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _0721_ (.A(_0331_),
    .B(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0722_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(\uut.in1[6] ),
    .A1(\uut.in2[6] ),
    .S(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _0724_ (.A(_0331_),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _0725_ (.A(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(\uut.in1[7] ),
    .A1(\uut.in2[7] ),
    .S(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(_0331_),
    .B(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0728_ (.A(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0340_));
 sky130_fd_sc_hd__a21oi_1 _0730_ (.A1(_0340_),
    .A2(net46),
    .B1(out_ready),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0341_));
 sky130_fd_sc_hd__nor2_1 _0731_ (.A(_0176_),
    .B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0054_));
 sky130_fd_sc_hd__or3b_1 _0732_ (.A(\count[1] ),
    .B(net1),
    .C_N(\count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__and3_1 _0733_ (.A(net46),
    .B(_0203_),
    .C(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__a31o_1 _0734_ (.A1(_0340_),
    .A2(_0307_),
    .A3(_0342_),
    .B1(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__a21oi_1 _0735_ (.A1(_0340_),
    .A2(_0342_),
    .B1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0056_));
 sky130_fd_sc_hd__and2_1 _0736_ (.A(_0331_),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _0738_ (.A(_0331_),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _0740_ (.A(_0331_),
    .B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _0741_ (.A(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _0742_ (.A(_0331_),
    .B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _0744_ (.A(_0331_),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _0745_ (.A(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _0746_ (.A(_0331_),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__clkbuf_2 _0748_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__and2_1 _0749_ (.A(_0350_),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0750_ (.A(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _0751_ (.A(_0350_),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _0752_ (.A(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__and2_1 _0753_ (.A(_0350_),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _0754_ (.A(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _0755_ (.A(_0350_),
    .B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0756_ (.A(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__and2_1 _0757_ (.A(_0350_),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0758_ (.A(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _0759_ (.A(_0350_),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0760_ (.A(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _0761_ (.A(_0350_),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _0762_ (.A(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _0763_ (.A(_0350_),
    .B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_1 _0764_ (.A(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _0765_ (.A(_0350_),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0766_ (.A(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _0767_ (.A(_0350_),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _0768_ (.A(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__buf_2 _0769_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _0770_ (.A(_0361_),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0771_ (.A(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _0772_ (.A(_0361_),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0773_ (.A(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _0774_ (.A(_0361_),
    .B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _0775_ (.A(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _0776_ (.A(_0361_),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0777_ (.A(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _0778_ (.A(_0361_),
    .B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0779_ (.A(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _0780_ (.A(_0361_),
    .B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _0781_ (.A(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _0782_ (.A(_0361_),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _0783_ (.A(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _0784_ (.A(_0361_),
    .B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0785_ (.A(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _0786_ (.A(_0361_),
    .B(\uut.mod_inv.inv_out1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0787_ (.A(_0370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _0788_ (.A(_0361_),
    .B(\uut.mod_inv.inv_out1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0789_ (.A(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_4 _0790_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__and2_1 _0791_ (.A(_0372_),
    .B(\uut.mod_inv.inv_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0792_ (.A(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _0793_ (.A(_0372_),
    .B(\uut.mod_inv.inv_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0794_ (.A(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__a21oi_1 _0795_ (.A1(\uut.R1[4] ),
    .A2(\uut.mod_inv.inv_out2[0] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0375_));
 sky130_fd_sc_hd__o21a_1 _0796_ (.A1(net93),
    .A2(\uut.mod_inv.inv_out2[0] ),
    .B1(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__a21oi_1 _0797_ (.A1(\uut.R1[5] ),
    .A2(\uut.mod_inv.inv_out2[1] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0376_));
 sky130_fd_sc_hd__o21a_1 _0798_ (.A1(\uut.R1[5] ),
    .A2(\uut.mod_inv.inv_out2[1] ),
    .B1(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__a21oi_1 _0799_ (.A1(\uut.R1[6] ),
    .A2(\uut.mod_inv.inv_out2[2] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0377_));
 sky130_fd_sc_hd__o21a_1 _0800_ (.A1(net81),
    .A2(\uut.mod_inv.inv_out2[2] ),
    .B1(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__a21oi_1 _0801_ (.A1(\uut.R1[7] ),
    .A2(\uut.mod_inv.inv_out2[3] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0378_));
 sky130_fd_sc_hd__o21a_1 _0802_ (.A1(net90),
    .A2(\uut.mod_inv.inv_out2[3] ),
    .B1(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__a21oi_1 _0803_ (.A1(\uut.R1[0] ),
    .A2(\uut.mod_inv.inv_out3[0] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0379_));
 sky130_fd_sc_hd__o21a_1 _0804_ (.A1(\uut.R1[0] ),
    .A2(\uut.mod_inv.inv_out3[0] ),
    .B1(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_1 _0805_ (.A1(\uut.R1[1] ),
    .A2(\uut.mod_inv.inv_out3[1] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0380_));
 sky130_fd_sc_hd__o21a_1 _0806_ (.A1(net80),
    .A2(\uut.mod_inv.inv_out3[1] ),
    .B1(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0090_));
 sky130_fd_sc_hd__a21oi_1 _0807_ (.A1(\uut.R1[2] ),
    .A2(\uut.mod_inv.inv_out3[2] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0381_));
 sky130_fd_sc_hd__o21a_1 _0808_ (.A1(net78),
    .A2(\uut.mod_inv.inv_out3[2] ),
    .B1(_0381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_1 _0809_ (.A1(\uut.R1[3] ),
    .A2(\uut.mod_inv.inv_out3[3] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0382_));
 sky130_fd_sc_hd__o21a_1 _0810_ (.A1(\uut.R1[3] ),
    .A2(\uut.mod_inv.inv_out3[3] ),
    .B1(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _0811_ (.A(_0372_),
    .B(\uut.mod_inv.inv_out4[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0812_ (.A(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _0813_ (.A(_0372_),
    .B(\uut.mod_inv.inv_out4[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _0814_ (.A(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _0815_ (.A(_0372_),
    .B(\uut.mod_inv.inv_out4[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _0816_ (.A(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _0817_ (.A(_0372_),
    .B(\uut.mod_inv.inv_out4[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _0818_ (.A(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__a21oi_1 _0819_ (.A1(\uut.R1[4] ),
    .A2(\uut.R1[0] ),
    .B1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0387_));
 sky130_fd_sc_hd__o21a_1 _0820_ (.A1(net93),
    .A2(\uut.R1[0] ),
    .B1(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_4 _0821_ (.A(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__a21oi_1 _0822_ (.A1(\uut.R1[5] ),
    .A2(\uut.R1[1] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0389_));
 sky130_fd_sc_hd__o21a_1 _0823_ (.A1(\uut.R1[5] ),
    .A2(net80),
    .B1(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__a21oi_1 _0824_ (.A1(\uut.R1[6] ),
    .A2(\uut.R1[2] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0390_));
 sky130_fd_sc_hd__o21a_1 _0825_ (.A1(\uut.R1[6] ),
    .A2(net78),
    .B1(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__a21oi_1 _0826_ (.A1(\uut.R1[7] ),
    .A2(\uut.R1[3] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0391_));
 sky130_fd_sc_hd__o21a_1 _0827_ (.A1(net90),
    .A2(\uut.R1[3] ),
    .B1(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _0828_ (.A(_0372_),
    .B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _0829_ (.A(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _0830_ (.A(_0372_),
    .B(\uut.sel_in_sh1.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0831_ (.A(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__and2_1 _0832_ (.A(_0372_),
    .B(\uut.sel_in_sh1.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _0833_ (.A(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _0834_ (.A(_0372_),
    .B(\uut.sel_in_sh1.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _0835_ (.A(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_2 _0836_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _0837_ (.A(_0396_),
    .B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _0838_ (.A(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__and2_1 _0839_ (.A(_0396_),
    .B(\uut.sel_in_sh2.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _0840_ (.A(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__and2_1 _0841_ (.A(_0396_),
    .B(\uut.sel_in_sh2.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _0842_ (.A(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__and2_1 _0843_ (.A(_0396_),
    .B(\uut.sel_in_sh2.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _0844_ (.A(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__and2_1 _0845_ (.A(_0396_),
    .B(\uut.sel_in_sh3.m4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0846_ (.A(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__and2_1 _0847_ (.A(_0396_),
    .B(\uut.sel_in_sh3.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0110_));
 sky130_fd_sc_hd__and2_1 _0849_ (.A(_0396_),
    .B(\uut.sel_in_sh3.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _0850_ (.A(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__and2_1 _0851_ (.A(_0396_),
    .B(\uut.sel_in_sh3.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _0852_ (.A(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0112_));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(_0396_),
    .B(\uut.sel_in_sh1.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0854_ (.A(_0405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0113_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(_0176_),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0114_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(\uut.in1[0] ),
    .B(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _0857_ (.A(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _0858_ (.A(_0396_),
    .B(\uut.sel_in_sh1.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0859_ (.A(_0407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_2 _0860_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0408_));
 sky130_fd_sc_hd__and2_1 _0861_ (.A(_0408_),
    .B(\uut.sel_in_sh2.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _0862_ (.A(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__nor2_1 _0863_ (.A(_0176_),
    .B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0118_));
 sky130_fd_sc_hd__and2_1 _0864_ (.A(_0408_),
    .B(\uut.sel_in_sh2.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _0865_ (.A(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0120_));
 sky130_fd_sc_hd__and2_1 _0866_ (.A(_0408_),
    .B(\uut.sel_in_sh3.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0867_ (.A(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _0868_ (.A(_0176_),
    .B(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0122_));
 sky130_fd_sc_hd__and2_1 _0869_ (.A(_0408_),
    .B(\uut.sel_in_sh3.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _0870_ (.A(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(_0408_),
    .B(\uut.mod_inv.sq_scl_out1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _0872_ (.A(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _0873_ (.A(_0408_),
    .B(\uut.mod_inv.sq_scl_out1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0126_));
 sky130_fd_sc_hd__and2_1 _0875_ (.A(_0408_),
    .B(\uut.mod_inv.sq_scl_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0876_ (.A(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(_0408_),
    .B(\uut.mod_inv.sq_scl_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _0878_ (.A(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__and2_1 _0879_ (.A(_0408_),
    .B(\uut.mod_inv.sq_scl_out2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _0880_ (.A(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__and2_1 _0881_ (.A(_0408_),
    .B(\uut.mod_inv.sq_scl_out2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _0882_ (.A(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _0883_ (.A(_0203_),
    .B(\uut.mod_inv.sq_scl_out2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _0884_ (.A(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(_0203_),
    .B(\uut.mod_inv.sq_scl_out2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _0886_ (.A(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0132_));
 sky130_fd_sc_hd__and2_1 _0887_ (.A(_0203_),
    .B(\uut.mod_inv.mod_mul1_out1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _0888_ (.A(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _0889_ (.A(_0203_),
    .B(\uut.mod_inv.mod_mul1_out1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _0890_ (.A(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _0891_ (.A(_0203_),
    .B(\uut.mod_inv.mod_mul1_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0892_ (.A(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _0893_ (.A(_0203_),
    .B(\uut.mod_inv.mod_mul1_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _0894_ (.A(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__a21oi_1 _0895_ (.A1(\uut.R0[4] ),
    .A2(\uut.mod_inv.mod_mul1_out2[0] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0425_));
 sky130_fd_sc_hd__o21a_1 _0896_ (.A1(net91),
    .A2(\uut.mod_inv.mod_mul1_out2[0] ),
    .B1(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0137_));
 sky130_fd_sc_hd__a21oi_1 _0897_ (.A1(\uut.R0[5] ),
    .A2(\uut.mod_inv.mod_mul1_out2[1] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0426_));
 sky130_fd_sc_hd__o21a_1 _0898_ (.A1(net84),
    .A2(\uut.mod_inv.mod_mul1_out2[1] ),
    .B1(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__a21oi_1 _0899_ (.A1(\uut.R0[6] ),
    .A2(\uut.mod_inv.mod_mul1_out2[2] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0427_));
 sky130_fd_sc_hd__o21a_1 _0900_ (.A1(net88),
    .A2(\uut.mod_inv.mod_mul1_out2[2] ),
    .B1(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__a21oi_1 _0901_ (.A1(net82),
    .A2(\uut.mod_inv.mod_mul1_out2[3] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0428_));
 sky130_fd_sc_hd__o21a_1 _0902_ (.A1(net82),
    .A2(\uut.mod_inv.mod_mul1_out2[3] ),
    .B1(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__a21oi_1 _0903_ (.A1(net72),
    .A2(\uut.mod_inv.mod_mul1_out3[0] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0429_));
 sky130_fd_sc_hd__o21a_1 _0904_ (.A1(net72),
    .A2(\uut.mod_inv.mod_mul1_out3[0] ),
    .B1(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__a21oi_1 _0905_ (.A1(net76),
    .A2(\uut.mod_inv.mod_mul1_out3[1] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0430_));
 sky130_fd_sc_hd__o21a_1 _0906_ (.A1(net76),
    .A2(\uut.mod_inv.mod_mul1_out3[1] ),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__a21oi_1 _0907_ (.A1(net87),
    .A2(\uut.mod_inv.mod_mul1_out3[2] ),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0431_));
 sky130_fd_sc_hd__o21a_1 _0908_ (.A1(net85),
    .A2(\uut.mod_inv.mod_mul1_out3[2] ),
    .B1(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__a21oi_1 _0909_ (.A1(net74),
    .A2(\uut.mod_inv.mod_mul1_out3[3] ),
    .B1(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0432_));
 sky130_fd_sc_hd__o21a_1 _0910_ (.A1(net74),
    .A2(\uut.mod_inv.mod_mul1_out3[3] ),
    .B1(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__dfxtp_1 _0911_ (.CLK(clknet_4_4_0_clk),
    .D(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0912_ (.CLK(clknet_4_4_0_clk),
    .D(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0913_ (.CLK(clknet_4_7_0_clk),
    .D(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0914_ (.CLK(clknet_4_4_0_clk),
    .D(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0915_ (.CLK(clknet_4_10_0_clk),
    .D(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_4 _0916_ (.CLK(clknet_4_10_0_clk),
    .D(_0005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_4 _0917_ (.CLK(clknet_4_10_0_clk),
    .D(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_4 _0918_ (.CLK(clknet_4_10_0_clk),
    .D(_0007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _0919_ (.CLK(clknet_4_10_0_clk),
    .D(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_4 _0920_ (.CLK(clknet_4_10_0_clk),
    .D(_0009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _0921_ (.CLK(clknet_4_10_0_clk),
    .D(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_4 _0922_ (.CLK(clknet_4_10_0_clk),
    .D(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfxtp_1 _0923_ (.CLK(clknet_4_11_0_clk),
    .D(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_count[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0924_ (.CLK(clknet_4_11_0_clk),
    .D(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_count[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0925_ (.CLK(clknet_4_11_0_clk),
    .D(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0926_ (.CLK(clknet_4_11_0_clk),
    .D(_0015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0927_ (.CLK(clknet_4_11_0_clk),
    .D(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0928_ (.CLK(clknet_4_11_0_clk),
    .D(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0929_ (.CLK(clknet_4_9_0_clk),
    .D(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0930_ (.CLK(clknet_4_11_0_clk),
    .D(_0019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0931_ (.CLK(clknet_4_11_0_clk),
    .D(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0932_ (.CLK(clknet_4_13_0_clk),
    .D(_0021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0933_ (.CLK(clknet_4_13_0_clk),
    .D(_0022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0934_ (.CLK(clknet_4_13_0_clk),
    .D(_0023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0935_ (.CLK(clknet_4_13_0_clk),
    .D(_0024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0936_ (.CLK(clknet_4_12_0_clk),
    .D(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0937_ (.CLK(clknet_4_13_0_clk),
    .D(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_4_13_0_clk),
    .D(_0027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_4_12_0_clk),
    .D(_0028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0940_ (.CLK(clknet_4_7_0_clk),
    .D(_0029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.R0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _0941_ (.CLK(clknet_4_13_0_clk),
    .D(_0030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0942_ (.CLK(clknet_4_7_0_clk),
    .D(_0031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0943_ (.CLK(clknet_4_6_0_clk),
    .D(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0944_ (.CLK(clknet_4_7_0_clk),
    .D(_0033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0945_ (.CLK(clknet_4_4_0_clk),
    .D(_0034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[4] ));
 sky130_fd_sc_hd__dfxtp_4 _0946_ (.CLK(clknet_4_7_0_clk),
    .D(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0947_ (.CLK(clknet_4_6_0_clk),
    .D(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0948_ (.CLK(clknet_4_6_0_clk),
    .D(_0037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_4_9_0_clk),
    .D(_0038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0950_ (.CLK(clknet_4_6_0_clk),
    .D(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0951_ (.CLK(clknet_4_3_0_clk),
    .D(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0952_ (.CLK(clknet_4_6_0_clk),
    .D(_0041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0953_ (.CLK(clknet_4_1_0_clk),
    .D(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _0954_ (.CLK(clknet_4_2_0_clk),
    .D(_0043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0955_ (.CLK(clknet_4_1_0_clk),
    .D(_0044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0956_ (.CLK(clknet_4_3_0_clk),
    .D(_0045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in2[7] ));
 sky130_fd_sc_hd__dfxtp_4 _0957_ (.CLK(clknet_4_9_0_clk),
    .D(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0958_ (.CLK(clknet_4_1_0_clk),
    .D(_0047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0959_ (.CLK(clknet_4_1_0_clk),
    .D(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_4_1_0_clk),
    .D(_0049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0961_ (.CLK(clknet_4_1_0_clk),
    .D(_0050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_4_1_0_clk),
    .D(_0051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _0963_ (.CLK(clknet_4_1_0_clk),
    .D(_0052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _0964_ (.CLK(clknet_4_2_0_clk),
    .D(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.in1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_4_11_0_clk),
    .D(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(out_ready));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_4_11_0_clk),
    .D(_0055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_4_11_0_clk),
    .D(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0968_ (.CLK(clknet_4_1_0_clk),
    .D(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_4_0_0_clk),
    .D(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_4_1_0_clk),
    .D(_0059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_4_0_0_clk),
    .D(_0060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_1[3] ));
 sky130_fd_sc_hd__dfxtp_4 _0972_ (.CLK(clknet_4_0_0_clk),
    .D(_0061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0973_ (.CLK(clknet_4_0_0_clk),
    .D(_0062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0974_ (.CLK(clknet_4_2_0_clk),
    .D(_0063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_1[2] ));
 sky130_fd_sc_hd__dfxtp_4 _0975_ (.CLK(clknet_4_2_0_clk),
    .D(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0976_ (.CLK(clknet_4_3_0_clk),
    .D(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0977_ (.CLK(clknet_4_2_0_clk),
    .D(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0978_ (.CLK(clknet_4_2_0_clk),
    .D(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0979_ (.CLK(clknet_4_2_0_clk),
    .D(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_4_3_0_clk),
    .D(_0069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_4_3_0_clk),
    .D(_0070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_4_3_0_clk),
    .D(_0071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_4_3_0_clk),
    .D(_0072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_1_2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0984_ (.CLK(clknet_4_3_0_clk),
    .D(_0073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0985_ (.CLK(clknet_4_3_0_clk),
    .D(_0074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0986_ (.CLK(clknet_4_8_0_clk),
    .D(_0075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_2[2] ));
 sky130_fd_sc_hd__dfxtp_4 _0987_ (.CLK(clknet_4_12_0_clk),
    .D(_0076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_1_2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0988_ (.CLK(clknet_4_6_0_clk),
    .D(_0077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _0989_ (.CLK(clknet_4_6_0_clk),
    .D(_0078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0990_ (.CLK(clknet_4_8_0_clk),
    .D(_0079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0991_ (.CLK(clknet_4_12_0_clk),
    .D(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_1_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_4_8_0_clk),
    .D(_0081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out1_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_4_8_0_clk),
    .D(_0082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out1_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_4_9_0_clk),
    .D(_0083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out1_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_4_15_0_clk),
    .D(_0084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out1_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_4_9_0_clk),
    .D(_0085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out2_xor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_4_9_0_clk),
    .D(_0086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out2_xor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_4_9_0_clk),
    .D(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out2_xor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_15_0_clk),
    .D(_0088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out2_xor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_12_0_clk),
    .D(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out3_xor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_12_0_clk),
    .D(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out3_xor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_4_12_0_clk),
    .D(_0091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out3_xor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_4_14_0_clk),
    .D(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out3_xor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_14_0_clk),
    .D(_0093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out4_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_4_15_0_clk),
    .D(_0094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out4_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_14_0_clk),
    .D(_0095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out4_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_4_8_0_clk),
    .D(_0096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_out4_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_4_15_0_clk),
    .D(_0097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_4_15_0_clk),
    .D(_0098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_4_14_0_clk),
    .D(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_4_14_0_clk),
    .D(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.random_xor_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_4_0_0_clk),
    .D(_0101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_4_0_0_clk),
    .D(_0102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_4_0_0_clk),
    .D(_0103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_4_0_0_clk),
    .D(_0104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_4_0_0_clk),
    .D(_0105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_4_0_0_clk),
    .D(_0106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_4_0_0_clk),
    .D(_0107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(clknet_4_0_0_clk),
    .D(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_4_2_0_clk),
    .D(_0109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_4_2_0_clk),
    .D(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_4_0_0_clk),
    .D(_0111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_4_0_0_clk),
    .D(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_4_2_0_clk),
    .D(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(clknet_4_3_0_clk),
    .D(_0114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_4_3_0_clk),
    .D(_0115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_4_3_0_clk),
    .D(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh1_reg_0_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_4_6_0_clk),
    .D(_0117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(clknet_4_3_0_clk),
    .D(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_4_8_0_clk),
    .D(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_4_6_0_clk),
    .D(_0120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh2_reg_0_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_4_6_0_clk),
    .D(_0121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_4_3_0_clk),
    .D(_0122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_4_8_0_clk),
    .D(_0123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_4_6_0_clk),
    .D(_0124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sh3_reg_0_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_4_5_0_clk),
    .D(_0125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_4_5_0_clk),
    .D(_0126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_4_5_0_clk),
    .D(_0127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1039_ (.CLK(clknet_4_5_0_clk),
    .D(_0128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_4_5_0_clk),
    .D(_0129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sq_scl_out2_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_4_4_0_clk),
    .D(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sq_scl_out2_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_4_7_0_clk),
    .D(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sq_scl_out2_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_4_5_0_clk),
    .D(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.sq_scl_out2_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_4_5_0_clk),
    .D(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out1_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_4_5_0_clk),
    .D(_0134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out1_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_4_5_0_clk),
    .D(_0135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out1_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_4_5_0_clk),
    .D(_0136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out1_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_4_4_0_clk),
    .D(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out2_xor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_4_5_0_clk),
    .D(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out2_xor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_4_5_0_clk),
    .D(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out2_xor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_4_5_0_clk),
    .D(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.mod_mul1_out2_xor[3] ));
 sky130_fd_sc_hd__dfxtp_4 _1052_ (.CLK(clknet_4_4_0_clk),
    .D(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in4[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1053_ (.CLK(clknet_4_4_0_clk),
    .D(_0142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in4[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1054_ (.CLK(clknet_4_4_0_clk),
    .D(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in4[2] ));
 sky130_fd_sc_hd__dfxtp_4 _1055_ (.CLK(clknet_4_4_0_clk),
    .D(_0144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uut.mod_inv.inv_in4[3] ));
 sky130_fd_sc_hd__clkbuf_4 _1071_ (.A(out_ready),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 fanout12 (.A(\uut.sel_in_sh2.m4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_4 fanout14 (.A(\uut.mod_inv.mul_in3[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 fanout15 (.A(\uut.mod_inv.mul_in3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(\uut.mod_inv.mul_in3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(\uut.mod_inv.mul_in3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 fanout18 (.A(\uut.mod_inv.mul_in3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(\uut.mod_inv.mul_in3[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(\uut.mod_inv.mul_in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout22 (.A(\uut.mod_inv.inv_out3_xor[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_4 fanout23 (.A(\uut.mod_inv.inv_out3_xor[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(\uut.mod_inv.inv_out3_xor[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(\uut.mod_inv.inv_out3_xor[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_4 fanout26 (.A(\uut.mod_inv.inv_out3_xor[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_8 fanout27 (.A(\uut.in2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(\uut.in3[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\uut.mod_inv.sh1_reg_0_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\uut.mod_inv.sh1_reg_0_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\uut.mod_inv.sh3_reg_0_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\uut.mod_inv.sh1_reg_0_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\uut.mod_inv.sh3_reg_0_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\uut.mod_inv.sh1_reg_0_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\uut.mod_inv.sh3_reg_0_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\uut.mod_inv.sh2_reg_0_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\uut.mod_inv.sh1_reg_0_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\uut.mod_inv.sh2_reg_0_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\uut.mod_inv.sh3_reg_0_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\uut.mod_inv.sh3_reg_0_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\uut.mod_inv.sh2_reg_0_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\uut.mod_inv.sh1_reg_0_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\uut.mod_inv.sh3_reg_0_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\uut.mod_inv.sh1_reg_0_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\uut.mod_inv.sh2_reg_0_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\uut.mod_inv.sh1_reg_0_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\uut.mod_inv.sh2_reg_0_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\uut.mod_inv.sh2_reg_0_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\uut.mod_inv.sh2_reg_0_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_1 hold29 (.A(\uut.R0[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_1 hold31 (.A(\uut.R0[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_1 hold33 (.A(\uut.R0[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__buf_1 hold35 (.A(\uut.R1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__buf_1 hold37 (.A(\uut.R1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\uut.R1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\uut.R0[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(out_ready),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\uut.R0[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\uut.R0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\uut.R0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\uut.R0[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\out_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\uut.R1[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\uut.R0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\uut.in2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\uut.R1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(uo_out[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\uut.mod_inv.sh3_reg_0_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\uut.mod_inv.sh2_reg_0_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\uut.mod_inv.sh3_reg_0_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap1 (.A(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__buf_4 max_cap11 (.A(\uut.sel_in_sh1.m4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_4 max_cap13 (.A(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_4 max_cap21 (.A(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__conb_1 tt_um_prg_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net29));
 sky130_fd_sc_hd__conb_1 tt_um_prg_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__conb_1 tt_um_prg_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__conb_1 tt_um_prg_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__conb_1 tt_um_prg_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net33));
 sky130_fd_sc_hd__conb_1 tt_um_prg_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_prg_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_prg_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net36));
 sky130_fd_sc_hd__conb_1 tt_um_prg_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net37));
 sky130_fd_sc_hd__conb_1 tt_um_prg_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net38));
 sky130_fd_sc_hd__conb_1 tt_um_prg_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net39));
 sky130_fd_sc_hd__conb_1 tt_um_prg_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net40));
 sky130_fd_sc_hd__conb_1 tt_um_prg_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net41));
 sky130_fd_sc_hd__conb_1 tt_um_prg_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net42));
 sky130_fd_sc_hd__conb_1 tt_um_prg_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net43));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_255_  (.A(\uut.mod_inv.inv_in3[0] ),
    .B(\uut.mod_inv.inv_in4[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_190_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.inv_mod/_256_  (.A(\uut.mod_inv.inv_mod/_190_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_191_ ));
 sky130_fd_sc_hd__inv_2 \uut.mod_inv.inv_mod/_257_  (.A(\uut.mod_inv.inv_in2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_192_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_258_  (.A(\uut.mod_inv.inv_in2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_193_ ));
 sky130_fd_sc_hd__clkbuf_8 \uut.mod_inv.inv_mod/_259_  (.A(\uut.mod_inv.inv_in3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_194_ ));
 sky130_fd_sc_hd__xor2_4 \uut.mod_inv.inv_mod/_260_  (.A(\uut.mod_inv.inv_mod/_194_ ),
    .B(\uut.mod_inv.inv_in4[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_195_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_261_  (.A(\uut.mod_inv.inv_mod/_193_ ),
    .B(\uut.mod_inv.inv_mod/_195_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_196_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_262_  (.A(\uut.mod_inv.inv_in2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_197_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.inv_mod/_263_  (.A(\uut.mod_inv.inv_in3[1] ),
    .B(\uut.mod_inv.inv_in4[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_198_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_264_  (.A(\uut.mod_inv.inv_mod/_197_ ),
    .B(\uut.mod_inv.inv_mod/_198_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_199_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_265_  (.A(\uut.mod_inv.inv_mod/_196_ ),
    .B(\uut.mod_inv.inv_mod/_199_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_200_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_266_  (.A0(\uut.mod_inv.inv_mod/_191_ ),
    .A1(\uut.mod_inv.inv_mod/_192_ ),
    .S(\uut.mod_inv.inv_mod/_200_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_201_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_267_  (.A(\uut.mod_inv.inv_in2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_202_ ));
 sky130_fd_sc_hd__xor2_4 \uut.mod_inv.inv_mod/_268_  (.A(\uut.mod_inv.inv_in3[3] ),
    .B(\uut.mod_inv.inv_in4[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_203_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_269_  (.A(\uut.mod_inv.inv_mod/_202_ ),
    .B(\uut.mod_inv.inv_mod/_203_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_204_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_270_  (.A0(\uut.mod_inv.inv_mod/_198_ ),
    .A1(\uut.mod_inv.inv_mod/_197_ ),
    .S(\uut.mod_inv.inv_mod/_204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_205_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_271_  (.A(\uut.mod_inv.inv_mod/_201_ ),
    .B(\uut.mod_inv.inv_mod/_205_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out1[3] ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_272_  (.A(\uut.mod_inv.inv_in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_206_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_273_  (.A(\uut.mod_inv.inv_mod/_206_ ),
    .B(\uut.mod_inv.inv_mod/_195_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_207_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_274_  (.A(\uut.mod_inv.inv_mod/_191_ ),
    .B(\uut.mod_inv.inv_mod/_207_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_208_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_275_  (.A(\uut.mod_inv.inv_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_209_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_276_  (.A(\uut.mod_inv.inv_mod/_206_ ),
    .B(\uut.mod_inv.inv_mod/_203_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_210_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_277_  (.A(\uut.mod_inv.inv_mod/_206_ ),
    .B(\uut.mod_inv.inv_mod/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_211_ ));
 sky130_fd_sc_hd__o22a_2 \uut.mod_inv.inv_mod/_278_  (.A1(\uut.mod_inv.inv_mod/_209_ ),
    .A2(\uut.mod_inv.inv_mod/_210_ ),
    .B1(\uut.mod_inv.inv_mod/_211_ ),
    .B2(\uut.mod_inv.inv_mod/_203_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_212_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_279_  (.A(\uut.mod_inv.inv_mod/_208_ ),
    .B(\uut.mod_inv.inv_mod/_212_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_213_ ));
 sky130_fd_sc_hd__buf_4 \uut.mod_inv.inv_mod/_280_  (.A(\uut.mod_inv.inv_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_214_ ));
 sky130_fd_sc_hd__and3b_1 \uut.mod_inv.inv_mod/_281_  (.A_N(\uut.mod_inv.inv_mod/_191_ ),
    .B(\uut.mod_inv.inv_mod/_206_ ),
    .C(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_215_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_282_  (.A(\uut.mod_inv.inv_in1[2] ),
    .B(\uut.mod_inv.inv_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_216_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_283_  (.A0(\uut.mod_inv.inv_in4[1] ),
    .A1(\uut.mod_inv.inv_in3[1] ),
    .S(\uut.mod_inv.inv_mod/_216_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_217_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_284_  (.A(\uut.mod_inv.inv_mod/_215_ ),
    .B(\uut.mod_inv.inv_mod/_217_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_218_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_285_  (.A(\uut.mod_inv.inv_mod/_214_ ),
    .B(\uut.mod_inv.inv_mod/_195_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_219_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_286_  (.A(\uut.mod_inv.inv_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_220_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_287_  (.A(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_221_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.inv_mod/_288_  (.A(\uut.mod_inv.inv_mod/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_222_ ));
 sky130_fd_sc_hd__and3b_1 \uut.mod_inv.inv_mod/_289_  (.A_N(\uut.mod_inv.inv_mod/_219_ ),
    .B(\uut.mod_inv.inv_mod/_221_ ),
    .C(\uut.mod_inv.inv_mod/_222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_223_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_290_  (.A(\uut.mod_inv.inv_mod/_218_ ),
    .B(\uut.mod_inv.inv_mod/_223_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_224_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_291_  (.A(\uut.mod_inv.inv_mod/_213_ ),
    .B(\uut.mod_inv.inv_mod/_224_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_225_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_292_  (.A(\uut.mod_inv.inv_mod/_220_ ),
    .B(\uut.mod_inv.inv_mod/_195_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_226_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_293_  (.A(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_227_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_294_  (.A(\uut.mod_inv.inv_mod/_227_ ),
    .B(\uut.mod_inv.inv_mod/_191_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_228_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_295_  (.A(\uut.mod_inv.inv_in3[1] ),
    .B(\uut.mod_inv.inv_in4[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_229_ ));
 sky130_fd_sc_hd__a21oi_1 \uut.mod_inv.inv_mod/_296_  (.A1(\uut.mod_inv.inv_mod/_226_ ),
    .A2(\uut.mod_inv.inv_mod/_228_ ),
    .B1(\uut.mod_inv.inv_mod/_229_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_230_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_297_  (.A1(\uut.mod_inv.inv_mod/_226_ ),
    .A2(\uut.mod_inv.inv_mod/_228_ ),
    .B1(\uut.mod_inv.inv_mod/_230_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_231_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_298_  (.A(\uut.mod_inv.inv_mod/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_232_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_299_  (.A(\uut.mod_inv.inv_mod/_232_ ),
    .B(\uut.mod_inv.inv_mod/_229_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_233_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_300_  (.A(\uut.mod_inv.inv_mod/_209_ ),
    .B(\uut.mod_inv.inv_mod/_198_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_234_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_301_  (.A(\uut.mod_inv.inv_mod/_227_ ),
    .B(\uut.mod_inv.inv_mod/_234_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_235_ ));
 sky130_fd_sc_hd__a21oi_1 \uut.mod_inv.inv_mod/_302_  (.A1(\uut.mod_inv.inv_mod/_227_ ),
    .A2(\uut.mod_inv.inv_mod/_233_ ),
    .B1(\uut.mod_inv.inv_mod/_235_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_236_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_303_  (.A(\uut.mod_inv.inv_in3[0] ),
    .B(\uut.mod_inv.inv_mod/_236_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_237_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_304_  (.A(\uut.mod_inv.inv_mod/_231_ ),
    .B(\uut.mod_inv.inv_mod/_237_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_238_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_305_  (.A(\uut.mod_inv.inv_mod/_225_ ),
    .B(\uut.mod_inv.inv_mod/_238_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out2[3] ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_306_  (.A(\uut.mod_inv.inv_in2[2] ),
    .B(\uut.mod_inv.inv_mod/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_239_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_307_  (.A(\uut.mod_inv.inv_in4[0] ),
    .B(\uut.mod_inv.inv_mod/_239_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_240_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_308_  (.A(\uut.mod_inv.inv_in4[1] ),
    .B(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_241_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_309_  (.A(\uut.mod_inv.inv_in2[2] ),
    .B(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_242_ ));
 sky130_fd_sc_hd__inv_2 \uut.mod_inv.inv_mod/_310_  (.A(\uut.mod_inv.inv_in2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_243_ ));
 sky130_fd_sc_hd__inv_2 \uut.mod_inv.inv_mod/_311_  (.A(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_244_ ));
 sky130_fd_sc_hd__o2bb2a_1 \uut.mod_inv.inv_mod/_312_  (.A1_N(\uut.mod_inv.inv_mod/_216_ ),
    .A2_N(\uut.mod_inv.inv_mod/_242_ ),
    .B1(\uut.mod_inv.inv_mod/_243_ ),
    .B2(\uut.mod_inv.inv_mod/_244_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_245_ ));
 sky130_fd_sc_hd__inv_2 \uut.mod_inv.inv_mod/_313_  (.A(\uut.mod_inv.inv_in2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_246_ ));
 sky130_fd_sc_hd__o211a_1 \uut.mod_inv.inv_mod/_314_  (.A1(\uut.mod_inv.inv_mod/_246_ ),
    .A2(\uut.mod_inv.inv_mod/_216_ ),
    .B1(\uut.mod_inv.inv_mod/_242_ ),
    .C1(\uut.mod_inv.inv_in4[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_247_ ));
 sky130_fd_sc_hd__a31o_1 \uut.mod_inv.inv_mod/_315_  (.A1(\uut.mod_inv.inv_mod/_197_ ),
    .A2(\uut.mod_inv.inv_mod/_241_ ),
    .A3(\uut.mod_inv.inv_mod/_245_ ),
    .B1(\uut.mod_inv.inv_mod/_247_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_248_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_316_  (.A(\uut.mod_inv.inv_mod/_240_ ),
    .B(\uut.mod_inv.inv_mod/_248_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_249_ ));
 sky130_fd_sc_hd__a21oi_1 \uut.mod_inv.inv_mod/_317_  (.A1(\uut.mod_inv.inv_mod/_241_ ),
    .A2(\uut.mod_inv.inv_mod/_239_ ),
    .B1(\uut.mod_inv.inv_mod/_192_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_250_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_318_  (.A1(\uut.mod_inv.inv_mod/_241_ ),
    .A2(\uut.mod_inv.inv_mod/_239_ ),
    .B1(\uut.mod_inv.inv_mod/_250_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_251_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_319_  (.A(\uut.mod_inv.inv_in2[3] ),
    .B(\uut.mod_inv.inv_in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_252_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_320_  (.A(\uut.mod_inv.inv_mod/_197_ ),
    .B(\uut.mod_inv.inv_in4[2] ),
    .C(\uut.mod_inv.inv_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_253_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_321_  (.A(\uut.mod_inv.inv_mod/_252_ ),
    .B(\uut.mod_inv.inv_mod/_253_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_254_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_322_  (.A(\uut.mod_inv.inv_in2[0] ),
    .B(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_000_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_323_  (.A(\uut.mod_inv.inv_mod/_246_ ),
    .B(\uut.mod_inv.inv_mod/_000_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_324_  (.A(\uut.mod_inv.inv_mod/_254_ ),
    .B(\uut.mod_inv.inv_mod/_001_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_325_  (.A(\uut.mod_inv.inv_mod/_251_ ),
    .B(\uut.mod_inv.inv_mod/_002_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_003_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_326_  (.A(\uut.mod_inv.inv_mod/_249_ ),
    .B(\uut.mod_inv.inv_mod/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_004_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.inv_mod/_327_  (.A(\uut.mod_inv.inv_in2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_005_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_328_  (.A(\uut.mod_inv.inv_mod/_005_ ),
    .B(\uut.mod_inv.inv_in4[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_006_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_329_  (.A(\uut.mod_inv.inv_mod/_005_ ),
    .B(\uut.mod_inv.inv_in4[2] ),
    .C(\uut.mod_inv.inv_mod/_222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_007_ ));
 sky130_fd_sc_hd__o211a_1 \uut.mod_inv.inv_mod/_330_  (.A1(\uut.mod_inv.inv_mod/_192_ ),
    .A2(\uut.mod_inv.inv_mod/_243_ ),
    .B1(\uut.mod_inv.inv_mod/_227_ ),
    .C1(\uut.mod_inv.inv_mod/_222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_008_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_331_  (.A1(\uut.mod_inv.inv_mod/_005_ ),
    .A2(\uut.mod_inv.inv_mod/_193_ ),
    .B1(\uut.mod_inv.inv_mod/_008_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_009_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_332_  (.A0(\uut.mod_inv.inv_mod/_006_ ),
    .A1(\uut.mod_inv.inv_mod/_007_ ),
    .S(\uut.mod_inv.inv_mod/_009_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_010_ ));
 sky130_fd_sc_hd__nand2_4 \uut.mod_inv.inv_mod/_333_  (.A(\uut.mod_inv.inv_mod/_197_ ),
    .B(\uut.mod_inv.inv_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_011_ ));
 sky130_fd_sc_hd__and2_1 \uut.mod_inv.inv_mod/_334_  (.A(\uut.mod_inv.inv_in2[1] ),
    .B(\uut.mod_inv.inv_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_012_ ));
 sky130_fd_sc_hd__clkbuf_2 \uut.mod_inv.inv_mod/_335_  (.A(\uut.mod_inv.inv_mod/_012_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_013_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_336_  (.A(\uut.mod_inv.inv_in4[0] ),
    .B(\uut.mod_inv.inv_mod/_013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_014_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_337_  (.A(\uut.mod_inv.inv_mod/_011_ ),
    .B(\uut.mod_inv.inv_mod/_014_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_015_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_338_  (.A(\uut.mod_inv.inv_mod/_010_ ),
    .B(\uut.mod_inv.inv_mod/_015_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_016_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_339_  (.A(\uut.mod_inv.inv_mod/_004_ ),
    .B(\uut.mod_inv.inv_mod/_016_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out3[3] ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_340_  (.A(\uut.mod_inv.inv_in3[1] ),
    .B(\uut.mod_inv.inv_mod/_193_ ),
    .C(\uut.mod_inv.inv_mod/_221_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_017_ ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_341_  (.A1(\uut.mod_inv.inv_mod/_005_ ),
    .A2(\uut.mod_inv.inv_mod/_194_ ),
    .B1_N(\uut.mod_inv.inv_mod/_222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_342_  (.A(\uut.mod_inv.inv_mod/_017_ ),
    .B(\uut.mod_inv.inv_mod/_018_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_019_ ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_343_  (.A1(\uut.mod_inv.inv_mod/_197_ ),
    .A2(\uut.mod_inv.inv_mod/_194_ ),
    .B1_N(\uut.mod_inv.inv_mod/_221_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_020_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_344_  (.A(\uut.mod_inv.inv_mod/_005_ ),
    .B(\uut.mod_inv.inv_in3[1] ),
    .C(\uut.mod_inv.inv_mod/_227_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_021_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_345_  (.A(\uut.mod_inv.inv_mod/_020_ ),
    .B(\uut.mod_inv.inv_mod/_021_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_022_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_346_  (.A(\uut.mod_inv.inv_mod/_019_ ),
    .B(\uut.mod_inv.inv_mod/_022_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_023_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_347_  (.A(\uut.mod_inv.inv_mod/_239_ ),
    .B(\uut.mod_inv.inv_mod/_013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_024_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_348_  (.A(\uut.mod_inv.inv_in3[0] ),
    .B(\uut.mod_inv.inv_mod/_024_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_025_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_349_  (.A(\uut.mod_inv.inv_mod/_023_ ),
    .B(\uut.mod_inv.inv_mod/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out4[3] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_350_  (.A(\uut.mod_inv.inv_in2[0] ),
    .B(\uut.mod_inv.inv_mod/_191_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_026_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_351_  (.A(\uut.mod_inv.inv_mod/_199_ ),
    .B(\uut.mod_inv.inv_mod/_204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_027_ ));
 sky130_fd_sc_hd__o21a_1 \uut.mod_inv.inv_mod/_352_  (.A1(\uut.mod_inv.inv_mod/_196_ ),
    .A2(\uut.mod_inv.inv_mod/_026_ ),
    .B1(\uut.mod_inv.inv_mod/_027_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_028_ ));
 sky130_fd_sc_hd__o2bb2a_1 \uut.mod_inv.inv_mod/_353_  (.A1_N(\uut.mod_inv.inv_mod/_200_ ),
    .A2_N(\uut.mod_inv.inv_mod/_028_ ),
    .B1(\uut.mod_inv.inv_mod/_026_ ),
    .B2(\uut.mod_inv.inv_mod/_027_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_029_ ));
 sky130_fd_sc_hd__o21a_1 \uut.mod_inv.inv_mod/_354_  (.A1(\uut.mod_inv.inv_mod/_200_ ),
    .A2(\uut.mod_inv.inv_mod/_028_ ),
    .B1(\uut.mod_inv.inv_mod/_029_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_030_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_355_  (.A(\uut.mod_inv.inv_mod/_192_ ),
    .B(\uut.mod_inv.inv_mod/_030_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out1[2] ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_356_  (.A(\uut.mod_inv.inv_mod/_220_ ),
    .B(\uut.mod_inv.inv_mod/_203_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_031_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_357_  (.A(\uut.mod_inv.inv_mod/_209_ ),
    .B(\uut.mod_inv.inv_mod/_191_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_032_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_358_  (.A(\uut.mod_inv.inv_mod/_031_ ),
    .B(\uut.mod_inv.inv_mod/_032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_033_ ));
 sky130_fd_sc_hd__a211o_1 \uut.mod_inv.inv_mod/_359_  (.A1(\uut.mod_inv.inv_mod/_031_ ),
    .A2(\uut.mod_inv.inv_mod/_032_ ),
    .B1(\uut.mod_inv.inv_mod/_033_ ),
    .C1(\uut.mod_inv.inv_mod/_229_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_034_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_360_  (.A(\uut.mod_inv.inv_mod/_194_ ),
    .B(\uut.mod_inv.inv_in4[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_035_ ));
 sky130_fd_sc_hd__nand2_2 \uut.mod_inv.inv_mod/_361_  (.A(\uut.mod_inv.inv_in1[3] ),
    .B(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_036_ ));
 sky130_fd_sc_hd__o22a_1 \uut.mod_inv.inv_mod/_362_  (.A1(\uut.mod_inv.inv_mod/_221_ ),
    .A2(\uut.mod_inv.inv_mod/_035_ ),
    .B1(\uut.mod_inv.inv_mod/_229_ ),
    .B2(\uut.mod_inv.inv_mod/_036_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_363_  (.A(\uut.mod_inv.inv_mod/_034_ ),
    .B(\uut.mod_inv.inv_mod/_037_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_038_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_364_  (.A0(\uut.mod_inv.inv_in4[0] ),
    .A1(\uut.mod_inv.inv_in3[0] ),
    .S(\uut.mod_inv.inv_mod/_211_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_039_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_365_  (.A(\uut.mod_inv.inv_mod/_191_ ),
    .B(\uut.mod_inv.inv_mod/_210_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_040_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_366_  (.A0(\uut.mod_inv.inv_mod/_191_ ),
    .A1(\uut.mod_inv.inv_mod/_220_ ),
    .S(\uut.mod_inv.inv_mod/_210_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_041_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_367_  (.A(\uut.mod_inv.inv_mod/_244_ ),
    .B(\uut.mod_inv.inv_mod/_221_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_042_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_368_  (.A0(\uut.mod_inv.inv_mod/_040_ ),
    .A1(\uut.mod_inv.inv_mod/_041_ ),
    .S(\uut.mod_inv.inv_mod/_042_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_043_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_369_  (.A(\uut.mod_inv.inv_mod/_039_ ),
    .B(\uut.mod_inv.inv_mod/_043_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_044_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_370_  (.A(\uut.mod_inv.inv_mod/_038_ ),
    .B(\uut.mod_inv.inv_mod/_044_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_045_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_371_  (.A0(\uut.mod_inv.inv_mod/_233_ ),
    .A1(\uut.mod_inv.inv_mod/_236_ ),
    .S(\uut.mod_inv.inv_mod/_228_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_046_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_372_  (.A(\uut.mod_inv.inv_mod/_244_ ),
    .B(\uut.mod_inv.inv_mod/_036_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_047_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_373_  (.A0(\uut.mod_inv.inv_mod/_035_ ),
    .A1(\uut.mod_inv.inv_mod/_047_ ),
    .S(\uut.mod_inv.inv_mod/_222_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_048_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_374_  (.A(\uut.mod_inv.inv_mod/_212_ ),
    .B(\uut.mod_inv.inv_mod/_048_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_375_  (.A(\uut.mod_inv.inv_mod/_046_ ),
    .B(\uut.mod_inv.inv_mod/_049_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_050_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_376_  (.A(\uut.mod_inv.inv_mod/_045_ ),
    .B(\uut.mod_inv.inv_mod/_050_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out2[2] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_377_  (.A(\uut.mod_inv.inv_in4[1] ),
    .B(\uut.mod_inv.inv_in2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_051_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_378_  (.A1(\uut.mod_inv.inv_mod/_243_ ),
    .A2(\uut.mod_inv.inv_mod/_051_ ),
    .B1(\uut.mod_inv.inv_mod/_221_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_052_ ));
 sky130_fd_sc_hd__a21o_1 \uut.mod_inv.inv_mod/_379_  (.A1(\uut.mod_inv.inv_mod/_243_ ),
    .A2(\uut.mod_inv.inv_mod/_051_ ),
    .B1(\uut.mod_inv.inv_mod/_052_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_053_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_380_  (.A(\uut.mod_inv.inv_in2[0] ),
    .B(\uut.mod_inv.inv_in4[3] ),
    .C(\uut.mod_inv.inv_mod/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_054_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_381_  (.A(\uut.mod_inv.inv_in4[0] ),
    .B(\uut.mod_inv.inv_mod/_011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_055_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_382_  (.A(\uut.mod_inv.inv_mod/_054_ ),
    .B(\uut.mod_inv.inv_mod/_055_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_056_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_383_  (.A(\uut.mod_inv.inv_mod/_053_ ),
    .B(\uut.mod_inv.inv_mod/_056_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_057_ ));
 sky130_fd_sc_hd__nand3_1 \uut.mod_inv.inv_mod/_384_  (.A(\uut.mod_inv.inv_mod/_005_ ),
    .B(\uut.mod_inv.inv_in4[1] ),
    .C(\uut.mod_inv.inv_mod/_232_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_058_ ));
 sky130_fd_sc_hd__a32o_1 \uut.mod_inv.inv_mod/_385_  (.A1(\uut.mod_inv.inv_in4[1] ),
    .A2(\uut.mod_inv.inv_mod/_227_ ),
    .A3(\uut.mod_inv.inv_mod/_232_ ),
    .B1(\uut.mod_inv.inv_mod/_000_ ),
    .B2(\uut.mod_inv.inv_mod/_058_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_059_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_386_  (.A(\uut.mod_inv.inv_mod/_057_ ),
    .B(\uut.mod_inv.inv_mod/_059_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_060_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_387_  (.A(\uut.mod_inv.inv_mod/_192_ ),
    .B(\uut.mod_inv.inv_mod/_252_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_061_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_388_  (.A0(\uut.mod_inv.inv_mod/_239_ ),
    .A1(\uut.mod_inv.inv_in2[2] ),
    .S(\uut.mod_inv.inv_mod/_061_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_062_ ));
 sky130_fd_sc_hd__inv_2 \uut.mod_inv.inv_mod/_389_  (.A(\uut.mod_inv.inv_in2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_063_ ));
 sky130_fd_sc_hd__a211o_1 \uut.mod_inv.inv_mod/_390_  (.A1(\uut.mod_inv.inv_mod/_192_ ),
    .A2(\uut.mod_inv.inv_mod/_063_ ),
    .B1(\uut.mod_inv.inv_mod/_211_ ),
    .C1(\uut.mod_inv.inv_mod/_061_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_064_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_391_  (.A(\uut.mod_inv.inv_mod/_062_ ),
    .B(\uut.mod_inv.inv_mod/_064_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_065_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_392_  (.A(\uut.mod_inv.inv_mod/_011_ ),
    .B(\uut.mod_inv.inv_mod/_065_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_066_ ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_393_  (.A1(\uut.mod_inv.inv_mod/_197_ ),
    .A2(\uut.mod_inv.inv_in4[3] ),
    .B1_N(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_067_ ));
 sky130_fd_sc_hd__and2_1 \uut.mod_inv.inv_mod/_394_  (.A(\uut.mod_inv.inv_in2[1] ),
    .B(\uut.mod_inv.inv_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_068_ ));
 sky130_fd_sc_hd__clkbuf_2 \uut.mod_inv.inv_mod/_395_  (.A(\uut.mod_inv.inv_mod/_068_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_069_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_396_  (.A1(\uut.mod_inv.inv_mod/_221_ ),
    .A2(\uut.mod_inv.inv_mod/_069_ ),
    .B1(\uut.mod_inv.inv_mod/_067_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_070_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_397_  (.A(\uut.mod_inv.inv_mod/_192_ ),
    .B(\uut.mod_inv.inv_mod/_069_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_071_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_398_  (.A0(\uut.mod_inv.inv_mod/_067_ ),
    .A1(\uut.mod_inv.inv_mod/_070_ ),
    .S(\uut.mod_inv.inv_mod/_071_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_072_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_399_  (.A(\uut.mod_inv.inv_mod/_202_ ),
    .B(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_073_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_400_  (.A1(\uut.mod_inv.inv_mod/_063_ ),
    .A2(\uut.mod_inv.inv_mod/_216_ ),
    .B1(\uut.mod_inv.inv_mod/_197_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_074_ ));
 sky130_fd_sc_hd__a21oi_1 \uut.mod_inv.inv_mod/_401_  (.A1(\uut.mod_inv.inv_mod/_244_ ),
    .A2(\uut.mod_inv.inv_mod/_073_ ),
    .B1(\uut.mod_inv.inv_mod/_074_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_075_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_402_  (.A(\uut.mod_inv.inv_in4[0] ),
    .B(\uut.mod_inv.inv_mod/_252_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_076_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_403_  (.A(\uut.mod_inv.inv_mod/_075_ ),
    .B(\uut.mod_inv.inv_mod/_076_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_404_  (.A(\uut.mod_inv.inv_mod/_072_ ),
    .B(\uut.mod_inv.inv_mod/_077_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_078_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_405_  (.A(\uut.mod_inv.inv_mod/_066_ ),
    .B(\uut.mod_inv.inv_mod/_078_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_079_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_406_  (.A(\uut.mod_inv.inv_mod/_060_ ),
    .B(\uut.mod_inv.inv_mod/_079_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out3[2] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_407_  (.A(\uut.mod_inv.inv_mod/_252_ ),
    .B(\uut.mod_inv.inv_mod/_069_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_080_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_408_  (.A(\uut.mod_inv.inv_in3[0] ),
    .B(\uut.mod_inv.inv_mod/_080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_081_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.inv_mod/_409_  (.A(\uut.mod_inv.inv_in3[1] ),
    .B(\uut.mod_inv.inv_in3[3] ),
    .C(\uut.mod_inv.inv_mod/_222_ ),
    .D(\uut.mod_inv.inv_mod/_232_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_082_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.inv_mod/_410_  (.A1(\uut.mod_inv.inv_in3[3] ),
    .A2(\uut.mod_inv.inv_mod/_222_ ),
    .B1(\uut.mod_inv.inv_mod/_232_ ),
    .B2(\uut.mod_inv.inv_in3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_083_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_411_  (.A(\uut.mod_inv.inv_mod/_082_ ),
    .B(\uut.mod_inv.inv_mod/_083_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_084_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_412_  (.A(\uut.mod_inv.inv_mod/_005_ ),
    .B(\uut.mod_inv.inv_mod/_084_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_085_ ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.inv_mod/_413_  (.A1(\uut.mod_inv.inv_mod/_197_ ),
    .A2(\uut.mod_inv.inv_in3[3] ),
    .B1(\uut.mod_inv.inv_mod/_202_ ),
    .B2(\uut.mod_inv.inv_in3[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_086_ ));
 sky130_fd_sc_hd__nand4_1 \uut.mod_inv.inv_mod/_414_  (.A(\uut.mod_inv.inv_in3[1] ),
    .B(\uut.mod_inv.inv_mod/_197_ ),
    .C(\uut.mod_inv.inv_in3[3] ),
    .D(\uut.mod_inv.inv_mod/_202_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_087_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_415_  (.A(\uut.mod_inv.inv_mod/_086_ ),
    .B(\uut.mod_inv.inv_mod/_087_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_088_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_416_  (.A(\uut.mod_inv.inv_mod/_221_ ),
    .B(\uut.mod_inv.inv_mod/_088_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_089_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_417_  (.A(\uut.mod_inv.inv_mod/_085_ ),
    .B(\uut.mod_inv.inv_mod/_089_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_090_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_418_  (.A(\uut.mod_inv.inv_mod/_081_ ),
    .B(\uut.mod_inv.inv_mod/_090_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out4[2] ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_419_  (.A(\uut.mod_inv.inv_mod/_204_ ),
    .B(\uut.mod_inv.inv_mod/_026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_091_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_420_  (.A0(\uut.mod_inv.inv_mod/_193_ ),
    .A1(\uut.mod_inv.inv_mod/_035_ ),
    .S(\uut.mod_inv.inv_mod/_091_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_092_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_421_  (.A(\uut.mod_inv.inv_mod/_232_ ),
    .B(\uut.mod_inv.inv_mod/_027_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_093_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_422_  (.A(\uut.mod_inv.inv_mod/_092_ ),
    .B(\uut.mod_inv.inv_mod/_093_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out1[1] ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_423_  (.A1(\uut.mod_inv.inv_mod/_191_ ),
    .A2(\uut.mod_inv.inv_mod/_203_ ),
    .B1_N(\uut.mod_inv.inv_mod/_036_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_094_ ));
 sky130_fd_sc_hd__o211a_1 \uut.mod_inv.inv_mod/_424_  (.A1(\uut.mod_inv.inv_mod/_031_ ),
    .A2(\uut.mod_inv.inv_mod/_032_ ),
    .B1(\uut.mod_inv.inv_mod/_094_ ),
    .C1(\uut.mod_inv.inv_mod/_227_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_095_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_425_  (.A(\uut.mod_inv.inv_mod/_202_ ),
    .B(\uut.mod_inv.inv_mod/_234_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_096_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_426_  (.A(\uut.mod_inv.inv_mod/_219_ ),
    .B(\uut.mod_inv.inv_mod/_032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_097_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_427_  (.A(\uut.mod_inv.inv_mod/_096_ ),
    .B(\uut.mod_inv.inv_mod/_097_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_098_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_428_  (.A(\uut.mod_inv.inv_mod/_095_ ),
    .B(\uut.mod_inv.inv_mod/_098_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_099_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_429_  (.A(\uut.mod_inv.inv_mod/_219_ ),
    .B(\uut.mod_inv.inv_mod/_031_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_100_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_430_  (.A(\uut.mod_inv.inv_mod/_194_ ),
    .B(\uut.mod_inv.inv_mod/_100_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_101_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_431_  (.A(\uut.mod_inv.inv_mod/_195_ ),
    .B(\uut.mod_inv.inv_mod/_036_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_102_ ));
 sky130_fd_sc_hd__a32o_1 \uut.mod_inv.inv_mod/_432_  (.A1(\uut.mod_inv.inv_mod/_221_ ),
    .A2(\uut.mod_inv.inv_mod/_035_ ),
    .A3(\uut.mod_inv.inv_mod/_191_ ),
    .B1(\uut.mod_inv.inv_mod/_032_ ),
    .B2(\uut.mod_inv.inv_mod/_102_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_103_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_433_  (.A(\uut.mod_inv.inv_mod/_212_ ),
    .B(\uut.mod_inv.inv_mod/_031_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_104_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_434_  (.A(\uut.mod_inv.inv_mod/_103_ ),
    .B(\uut.mod_inv.inv_mod/_104_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_105_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_435_  (.A(\uut.mod_inv.inv_mod/_101_ ),
    .B(\uut.mod_inv.inv_mod/_105_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_106_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_436_  (.A(\uut.mod_inv.inv_mod/_099_ ),
    .B(\uut.mod_inv.inv_mod/_106_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out2[1] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_437_  (.A(\uut.mod_inv.inv_in2[0] ),
    .B(\uut.mod_inv.inv_mod/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_107_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_438_  (.A(\uut.mod_inv.inv_mod/_202_ ),
    .B(\uut.mod_inv.inv_in4[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_108_ ));
 sky130_fd_sc_hd__o21a_1 \uut.mod_inv.inv_mod/_439_  (.A1(\uut.mod_inv.inv_mod/_107_ ),
    .A2(\uut.mod_inv.inv_mod/_108_ ),
    .B1(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_109_ ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_440_  (.A1(\uut.mod_inv.inv_mod/_107_ ),
    .A2(\uut.mod_inv.inv_mod/_108_ ),
    .B1_N(\uut.mod_inv.inv_mod/_109_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_110_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_441_  (.A(\uut.mod_inv.inv_in2[2] ),
    .B(\uut.mod_inv.inv_mod/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_111_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_442_  (.A(\uut.mod_inv.inv_mod/_192_ ),
    .B(\uut.mod_inv.inv_mod/_111_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_112_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_443_  (.A(\uut.mod_inv.inv_in2[0] ),
    .B(\uut.mod_inv.inv_in4[3] ),
    .C(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_113_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_444_  (.A0(\uut.mod_inv.inv_mod/_112_ ),
    .A1(\uut.mod_inv.inv_mod/_111_ ),
    .S(\uut.mod_inv.inv_mod/_113_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_114_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_445_  (.A(\uut.mod_inv.inv_mod/_110_ ),
    .B(\uut.mod_inv.inv_mod/_114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_115_ ));
 sky130_fd_sc_hd__and2_1 \uut.mod_inv.inv_mod/_446_  (.A(\uut.mod_inv.inv_mod/_202_ ),
    .B(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_116_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_447_  (.A(\uut.mod_inv.inv_in4[2] ),
    .B(\uut.mod_inv.inv_mod/_116_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_117_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_448_  (.A(\uut.mod_inv.inv_in4[2] ),
    .B(\uut.mod_inv.inv_mod/_202_ ),
    .C(\uut.mod_inv.inv_mod/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_118_ ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.inv_mod/_449_  (.A1(\uut.mod_inv.inv_mod/_252_ ),
    .A2(\uut.mod_inv.inv_mod/_117_ ),
    .B1(\uut.mod_inv.inv_mod/_118_ ),
    .B2(\uut.mod_inv.inv_mod/_221_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_119_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_450_  (.A(\uut.mod_inv.inv_mod/_116_ ),
    .B(\uut.mod_inv.inv_mod/_111_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_120_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_451_  (.A(\uut.mod_inv.inv_in2[2] ),
    .B(\uut.mod_inv.inv_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_121_ ));
 sky130_fd_sc_hd__o21a_1 \uut.mod_inv.inv_mod/_452_  (.A1(\uut.mod_inv.inv_in4[0] ),
    .A2(\uut.mod_inv.inv_mod/_111_ ),
    .B1(\uut.mod_inv.inv_mod/_121_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_122_ ));
 sky130_fd_sc_hd__o2bb2a_1 \uut.mod_inv.inv_mod/_453_  (.A1_N(\uut.mod_inv.inv_in4[0] ),
    .A2_N(\uut.mod_inv.inv_mod/_120_ ),
    .B1(\uut.mod_inv.inv_mod/_122_ ),
    .B2(\uut.mod_inv.inv_mod/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_123_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_454_  (.A(\uut.mod_inv.inv_mod/_119_ ),
    .B(\uut.mod_inv.inv_mod/_123_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_124_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_455_  (.A(\uut.mod_inv.inv_mod/_115_ ),
    .B(\uut.mod_inv.inv_mod/_124_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_125_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_456_  (.A(\uut.mod_inv.inv_mod/_063_ ),
    .B(\uut.mod_inv.inv_mod/_000_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_126_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_457_  (.A(\uut.mod_inv.inv_in3[3] ),
    .B(\uut.mod_inv.inv_mod/_126_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_127_ ));
 sky130_fd_sc_hd__a21oi_1 \uut.mod_inv.inv_mod/_458_  (.A1(\uut.mod_inv.inv_mod/_005_ ),
    .A2(\uut.mod_inv.inv_mod/_232_ ),
    .B1(\uut.mod_inv.inv_in4[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_128_ ));
 sky130_fd_sc_hd__and2_1 \uut.mod_inv.inv_mod/_459_  (.A(\uut.mod_inv.inv_mod/_246_ ),
    .B(\uut.mod_inv.inv_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_129_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_460_  (.A(\uut.mod_inv.inv_in4[3] ),
    .B(\uut.mod_inv.inv_mod/_129_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_130_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_461_  (.A0(\uut.mod_inv.inv_mod/_130_ ),
    .A1(\uut.mod_inv.inv_mod/_011_ ),
    .S(\uut.mod_inv.inv_mod/_242_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_131_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_462_  (.A(\uut.mod_inv.inv_mod/_128_ ),
    .B(\uut.mod_inv.inv_mod/_131_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_132_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_463_  (.A(\uut.mod_inv.inv_mod/_127_ ),
    .B(\uut.mod_inv.inv_mod/_132_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_133_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_464_  (.A(\uut.mod_inv.inv_mod/_125_ ),
    .B(\uut.mod_inv.inv_mod/_133_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out3[1] ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_465_  (.A1(\uut.mod_inv.inv_mod/_073_ ),
    .A2(\uut.mod_inv.inv_mod/_107_ ),
    .B1_N(\uut.mod_inv.inv_mod/_194_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_134_ ));
 sky130_fd_sc_hd__a31o_1 \uut.mod_inv.inv_mod/_466_  (.A1(\uut.mod_inv.inv_mod/_005_ ),
    .A2(\uut.mod_inv.inv_mod/_232_ ),
    .A3(\uut.mod_inv.inv_mod/_116_ ),
    .B1(\uut.mod_inv.inv_mod/_134_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_135_ ));
 sky130_fd_sc_hd__a21o_1 \uut.mod_inv.inv_mod/_467_  (.A1(\uut.mod_inv.inv_mod/_005_ ),
    .A2(\uut.mod_inv.inv_in3[3] ),
    .B1(\uut.mod_inv.inv_mod/_244_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_136_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_468_  (.A(\uut.mod_inv.inv_mod/_135_ ),
    .B(\uut.mod_inv.inv_mod/_136_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_137_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_469_  (.A0(\uut.mod_inv.inv_mod/_203_ ),
    .A1(\uut.mod_inv.inv_in4[3] ),
    .S(\uut.mod_inv.inv_mod/_242_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_138_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.inv_mod/_470_  (.A(\uut.mod_inv.inv_mod/_063_ ),
    .B(\uut.mod_inv.inv_mod/_244_ ),
    .C(\uut.mod_inv.inv_mod/_111_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_139_ ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.inv_mod/_471_  (.A1(\uut.mod_inv.inv_mod/_202_ ),
    .A2(\uut.mod_inv.inv_mod/_227_ ),
    .B1(\uut.mod_inv.inv_mod/_232_ ),
    .B2(\uut.mod_inv.inv_mod/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_140_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_472_  (.A(\uut.mod_inv.inv_in3[0] ),
    .B(\uut.mod_inv.inv_mod/_139_ ),
    .C(\uut.mod_inv.inv_mod/_140_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_141_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_473_  (.A(\uut.mod_inv.inv_mod/_138_ ),
    .B(\uut.mod_inv.inv_mod/_141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_142_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_474_  (.A(\uut.mod_inv.inv_mod/_137_ ),
    .B(\uut.mod_inv.inv_mod/_142_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out4[1] ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.inv_mod/_475_  (.A1(\uut.mod_inv.inv_mod/_200_ ),
    .A2(\uut.mod_inv.inv_mod/_204_ ),
    .B1_N(\uut.mod_inv.inv_mod/_028_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_143_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_476_  (.A0(\uut.mod_inv.inv_mod/_143_ ),
    .A1(\uut.mod_inv.inv_mod/_028_ ),
    .S(\uut.mod_inv.inv_mod/_091_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_144_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_477_  (.A(\uut.mod_inv.inv_mod/_243_ ),
    .B(\uut.mod_inv.inv_mod/_144_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out1[0] ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.inv_mod/_478_  (.A(\uut.mod_inv.inv_mod/_035_ ),
    .B(\uut.mod_inv.inv_mod/_210_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_145_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_479_  (.A(\uut.mod_inv.inv_mod/_216_ ),
    .B(\uut.mod_inv.inv_mod/_145_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_146_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.inv_mod/_480_  (.A(\uut.mod_inv.inv_mod/_244_ ),
    .B(\uut.mod_inv.inv_mod/_210_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_147_ ));
 sky130_fd_sc_hd__o22a_1 \uut.mod_inv.inv_mod/_481_  (.A1(\uut.mod_inv.inv_mod/_203_ ),
    .A2(\uut.mod_inv.inv_mod/_036_ ),
    .B1(\uut.mod_inv.inv_mod/_031_ ),
    .B2(\uut.mod_inv.inv_mod/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_148_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_482_  (.A(\uut.mod_inv.inv_mod/_147_ ),
    .B(\uut.mod_inv.inv_mod/_148_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_149_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_483_  (.A(\uut.mod_inv.inv_mod/_146_ ),
    .B(\uut.mod_inv.inv_mod/_149_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_150_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.inv_mod/_484_  (.A(\uut.mod_inv.inv_mod/_219_ ),
    .B(\uut.mod_inv.inv_mod/_234_ ),
    .C_N(\uut.mod_inv.inv_mod/_226_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_151_ ));
 sky130_fd_sc_hd__o21ai_1 \uut.mod_inv.inv_mod/_485_  (.A1(\uut.mod_inv.inv_mod/_226_ ),
    .A2(\uut.mod_inv.inv_mod/_235_ ),
    .B1(\uut.mod_inv.inv_mod/_151_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_152_ ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.inv_mod/_486_  (.A1(\uut.mod_inv.inv_mod/_198_ ),
    .A2(\uut.mod_inv.inv_mod/_203_ ),
    .B1_N(\uut.mod_inv.inv_mod/_211_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_153_ ));
 sky130_fd_sc_hd__o211a_1 \uut.mod_inv.inv_mod/_487_  (.A1(\uut.mod_inv.inv_mod/_210_ ),
    .A2(\uut.mod_inv.inv_mod/_234_ ),
    .B1(\uut.mod_inv.inv_mod/_153_ ),
    .C1(\uut.mod_inv.inv_mod/_227_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_154_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_488_  (.A(\uut.mod_inv.inv_mod/_152_ ),
    .B(\uut.mod_inv.inv_mod/_154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_155_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_489_  (.A(\uut.mod_inv.inv_mod/_150_ ),
    .B(\uut.mod_inv.inv_mod/_155_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_156_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_490_  (.A(\uut.mod_inv.inv_mod/_194_ ),
    .B(\uut.mod_inv.inv_mod/_212_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_157_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_491_  (.A(\uut.mod_inv.inv_mod/_232_ ),
    .B(\uut.mod_inv.inv_mod/_207_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_158_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_492_  (.A0(\uut.mod_inv.inv_mod/_209_ ),
    .A1(\uut.mod_inv.inv_mod/_214_ ),
    .S(\uut.mod_inv.inv_mod/_190_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_159_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_493_  (.A(\uut.mod_inv.inv_mod/_234_ ),
    .B(\uut.mod_inv.inv_mod/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_160_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_494_  (.A(\uut.mod_inv.inv_mod/_158_ ),
    .B(\uut.mod_inv.inv_mod/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_161_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_495_  (.A(\uut.mod_inv.inv_mod/_157_ ),
    .B(\uut.mod_inv.inv_mod/_161_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_162_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.inv_mod/_496_  (.A(\uut.mod_inv.inv_mod/_156_ ),
    .B(\uut.mod_inv.inv_mod/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out2[0] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_497_  (.A(\uut.mod_inv.inv_mod/_000_ ),
    .B(\uut.mod_inv.inv_mod/_011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_163_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_498_  (.A(\uut.mod_inv.inv_mod/_193_ ),
    .B(\uut.mod_inv.inv_in4[3] ),
    .C(\uut.mod_inv.inv_mod/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_164_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_499_  (.A(\uut.mod_inv.inv_in4[2] ),
    .B(\uut.mod_inv.inv_mod/_011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_165_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_500_  (.A(\uut.mod_inv.inv_mod/_164_ ),
    .B(\uut.mod_inv.inv_mod/_165_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_166_ ));
 sky130_fd_sc_hd__and3_1 \uut.mod_inv.inv_mod/_501_  (.A(\uut.mod_inv.inv_in4[1] ),
    .B(\uut.mod_inv.inv_mod/_193_ ),
    .C(\uut.mod_inv.inv_mod/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_167_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_502_  (.A(\uut.mod_inv.inv_mod/_116_ ),
    .B(\uut.mod_inv.inv_mod/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_168_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_503_  (.A(\uut.mod_inv.inv_mod/_166_ ),
    .B(\uut.mod_inv.inv_mod/_168_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_169_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_504_  (.A(\uut.mod_inv.inv_mod/_163_ ),
    .B(\uut.mod_inv.inv_mod/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_170_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_505_  (.A(\uut.mod_inv.inv_mod/_193_ ),
    .B(\uut.mod_inv.inv_mod/_069_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_171_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.inv_mod/_506_  (.A0(\uut.mod_inv.inv_in2[0] ),
    .A1(\uut.mod_inv.inv_mod/_107_ ),
    .S(\uut.mod_inv.inv_mod/_171_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_172_ ));
 sky130_fd_sc_hd__a21oi_1 \uut.mod_inv.inv_mod/_507_  (.A1(\uut.mod_inv.inv_mod/_222_ ),
    .A2(\uut.mod_inv.inv_mod/_013_ ),
    .B1(\uut.mod_inv.inv_mod/_063_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_173_ ));
 sky130_fd_sc_hd__o21a_1 \uut.mod_inv.inv_mod/_508_  (.A1(\uut.mod_inv.inv_mod/_222_ ),
    .A2(\uut.mod_inv.inv_mod/_013_ ),
    .B1(\uut.mod_inv.inv_mod/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_174_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_509_  (.A(\uut.mod_inv.inv_mod/_172_ ),
    .B(\uut.mod_inv.inv_mod/_174_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_175_ ));
 sky130_fd_sc_hd__a21o_1 \uut.mod_inv.inv_mod/_510_  (.A1(\uut.mod_inv.inv_mod/_206_ ),
    .A2(\uut.mod_inv.inv_in1[3] ),
    .B1(\uut.mod_inv.inv_mod/_220_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_176_ ));
 sky130_fd_sc_hd__o2111a_1 \uut.mod_inv.inv_mod/_511_  (.A1(\uut.mod_inv.inv_mod/_239_ ),
    .A2(\uut.mod_inv.inv_mod/_036_ ),
    .B1(\uut.mod_inv.inv_mod/_176_ ),
    .C1(\uut.mod_inv.inv_mod/_252_ ),
    .D1(\uut.mod_inv.inv_mod/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_177_ ));
 sky130_fd_sc_hd__a41o_1 \uut.mod_inv.inv_mod/_512_  (.A1(\uut.mod_inv.inv_mod/_202_ ),
    .A2(\uut.mod_inv.inv_mod/_222_ ),
    .A3(\uut.mod_inv.inv_mod/_242_ ),
    .A4(\uut.mod_inv.inv_mod/_121_ ),
    .B1(\uut.mod_inv.inv_mod/_177_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_178_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_513_  (.A(\uut.mod_inv.inv_in4[3] ),
    .B(\uut.mod_inv.inv_mod/_013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_179_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_514_  (.A(\uut.mod_inv.inv_mod/_118_ ),
    .B(\uut.mod_inv.inv_mod/_179_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_180_ ));
 sky130_fd_sc_hd__o21a_1 \uut.mod_inv.inv_mod/_515_  (.A1(\uut.mod_inv.inv_mod/_011_ ),
    .A2(\uut.mod_inv.inv_mod/_051_ ),
    .B1(\uut.mod_inv.inv_mod/_214_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_181_ ));
 sky130_fd_sc_hd__a21boi_1 \uut.mod_inv.inv_mod/_516_  (.A1(\uut.mod_inv.inv_mod/_011_ ),
    .A2(\uut.mod_inv.inv_mod/_051_ ),
    .B1_N(\uut.mod_inv.inv_mod/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_182_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_517_  (.A(\uut.mod_inv.inv_mod/_180_ ),
    .B(\uut.mod_inv.inv_mod/_182_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_183_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_518_  (.A(\uut.mod_inv.inv_mod/_178_ ),
    .B(\uut.mod_inv.inv_mod/_183_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_184_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_519_  (.A(\uut.mod_inv.inv_mod/_175_ ),
    .B(\uut.mod_inv.inv_mod/_184_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_185_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_520_  (.A(\uut.mod_inv.inv_mod/_170_ ),
    .B(\uut.mod_inv.inv_mod/_185_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out3[0] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_521_  (.A(\uut.mod_inv.inv_mod/_194_ ),
    .B(\uut.mod_inv.inv_mod/_080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_186_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_522_  (.A(\uut.mod_inv.inv_mod/_227_ ),
    .B(\uut.mod_inv.inv_mod/_088_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_187_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.inv_mod/_523_  (.A(\uut.mod_inv.inv_mod/_193_ ),
    .B(\uut.mod_inv.inv_mod/_084_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_mod/_188_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.inv_mod/_524_  (.A(\uut.mod_inv.inv_mod/_187_ ),
    .B(\uut.mod_inv.inv_mod/_188_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.inv_mod/_189_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.inv_mod/_525_  (.A(\uut.mod_inv.inv_mod/_186_ ),
    .B(\uut.mod_inv.inv_mod/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.inv_out4[0] ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul1/_221_  (.A(\uut.sel_in_sh3.m1.Q ),
    .B(\uut.sel_in_sh2.m1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_159_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul1/_222_  (.A(\uut.sel_in_sh3.m7.Q ),
    .B(\uut.sel_in_sh2.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_160_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul1/_223_  (.A(\uut.mod_inv.mod_mul1/_159_ ),
    .B(\uut.mod_inv.mod_mul1/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_161_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul1/_224_  (.A(\uut.sel_in_sh3.m6.Q ),
    .B(\uut.sel_in_sh2.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_162_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul1/_225_  (.A(net28),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_163_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_226_  (.A(\uut.mod_inv.mod_mul1/_162_ ),
    .B(\uut.mod_inv.mod_mul1/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_164_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_227_  (.A(\uut.mod_inv.mod_mul1/_161_ ),
    .B(\uut.mod_inv.mod_mul1/_164_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_165_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_228_  (.A(\uut.sel_in_sh3.m3.Q ),
    .B(\uut.sel_in_sh2.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_166_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul1/_229_  (.A(\uut.sel_in_sh3.m5.Q ),
    .B(\uut.sel_in_sh2.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_167_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_230_  (.A(\uut.mod_inv.mod_mul1/_166_ ),
    .B(\uut.mod_inv.mod_mul1/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_168_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_231_  (.A(\uut.sel_in_sh3.m5.Q ),
    .B(\uut.sel_in_sh2.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_169_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_232_  (.A(\uut.mod_inv.mod_mul1/_166_ ),
    .B(\uut.mod_inv.mod_mul1/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_170_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_233_  (.A0(\uut.mod_inv.mod_mul1/_168_ ),
    .A1(\uut.mod_inv.mod_mul1/_170_ ),
    .S(\uut.mod_inv.mod_mul1/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_171_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_234_  (.A(\uut.mod_inv.mod_mul1/_165_ ),
    .B(\uut.mod_inv.mod_mul1/_171_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_172_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_235_  (.A(\uut.sel_in_sh3.m0.Q ),
    .B(\uut.sel_in_sh2.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_173_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_236_  (.A(\uut.mod_inv.mod_mul1/_167_ ),
    .B(\uut.mod_inv.mod_mul1/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_174_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul1/_237_  (.A(\uut.mod_inv.mod_mul1/_169_ ),
    .B(\uut.mod_inv.mod_mul1/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_175_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_238_  (.A0(\uut.mod_inv.mod_mul1/_174_ ),
    .A1(\uut.mod_inv.mod_mul1/_175_ ),
    .S(\uut.mod_inv.mod_mul1/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_176_ ));
 sky130_fd_sc_hd__o22a_1 \uut.mod_inv.mod_mul1/_239_  (.A1(\uut.mod_inv.mod_mul1/_159_ ),
    .A2(\uut.mod_inv.mod_mul1/_162_ ),
    .B1(\uut.mod_inv.mod_mul1/_173_ ),
    .B2(\uut.mod_inv.mod_mul1/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_177_ ));
 sky130_fd_sc_hd__or4_1 \uut.mod_inv.mod_mul1/_240_  (.A(\uut.mod_inv.mod_mul1/_159_ ),
    .B(\uut.mod_inv.mod_mul1/_160_ ),
    .C(\uut.mod_inv.mod_mul1/_162_ ),
    .D(\uut.mod_inv.mod_mul1/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_178_ ));
 sky130_fd_sc_hd__nor2b_1 \uut.mod_inv.mod_mul1/_241_  (.A(\uut.mod_inv.mod_mul1/_177_ ),
    .B_N(\uut.mod_inv.mod_mul1/_178_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_179_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_242_  (.A(\uut.mod_inv.mod_mul1/_159_ ),
    .B(\uut.mod_inv.mod_mul1/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_180_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul1/_243_  (.A(\uut.sel_in_sh3.m4.Q ),
    .B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_181_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_244_  (.A0(\uut.mod_inv.mod_mul1/_167_ ),
    .A1(\uut.mod_inv.mod_mul1/_181_ ),
    .S(\uut.mod_inv.mod_mul1/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_182_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_245_  (.A(\uut.mod_inv.mod_mul1/_166_ ),
    .B(\uut.mod_inv.mod_mul1/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_183_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_246_  (.A0(\uut.mod_inv.mod_mul1/_180_ ),
    .A1(\uut.mod_inv.mod_mul1/_182_ ),
    .S(\uut.mod_inv.mod_mul1/_183_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_184_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_247_  (.A(\uut.mod_inv.mod_mul1/_179_ ),
    .B(\uut.mod_inv.mod_mul1/_184_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_185_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_248_  (.A(\uut.mod_inv.mod_mul1/_176_ ),
    .B(\uut.mod_inv.mod_mul1/_185_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_186_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_249_  (.A(\uut.mod_inv.mod_mul1/_172_ ),
    .B(\uut.mod_inv.mod_mul1/_186_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out1[3] ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_250_  (.A(\uut.sel_in_sh1.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_187_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_251_  (.A_N(\uut.sel_in_sh3.m0.Q ),
    .B(\uut.mod_inv.mod_mul1/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_188_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_252_  (.A(\uut.sel_in_sh1.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_189_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul1/_253_  (.A1(\uut.mod_inv.mod_mul1/_187_ ),
    .A2(\uut.mod_inv.mod_mul1/_189_ ),
    .B1_N(\uut.mod_inv.mod_mul1/_188_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_190_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_254_  (.A(\uut.sel_in_sh3.m7.Q ),
    .B_N(\uut.mod_inv.mod_mul1/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_191_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_255_  (.A0(\uut.mod_inv.mod_mul1/_188_ ),
    .A1(\uut.mod_inv.mod_mul1/_190_ ),
    .S(\uut.mod_inv.mod_mul1/_191_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_192_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_256_  (.A(\uut.sel_in_sh1.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_193_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_257_  (.A_N(\uut.sel_in_sh3.m1.Q ),
    .B(\uut.mod_inv.mod_mul1/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_194_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_258_  (.A0(\uut.sel_in_sh1.m1.Q ),
    .A1(\uut.sel_in_sh3.m1.Q ),
    .S(\uut.sel_in_sh1.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_195_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_259_  (.A(\uut.sel_in_sh3.m5.Q ),
    .B_N(\uut.sel_in_sh1.m1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_196_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_260_  (.A0(\uut.mod_inv.mod_mul1/_194_ ),
    .A1(\uut.mod_inv.mod_mul1/_195_ ),
    .S(\uut.mod_inv.mod_mul1/_196_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_197_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_261_  (.A_N(\uut.sel_in_sh3.m1.Q ),
    .B(\uut.sel_in_sh1.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_198_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_262_  (.A0(\uut.sel_in_sh1.m1.Q ),
    .A1(\uut.sel_in_sh3.m1.Q ),
    .S(\uut.sel_in_sh1.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_199_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_263_  (.A(\uut.sel_in_sh3.m7.Q ),
    .B_N(\uut.sel_in_sh1.m1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_200_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_264_  (.A0(\uut.mod_inv.mod_mul1/_198_ ),
    .A1(\uut.mod_inv.mod_mul1/_199_ ),
    .S(\uut.mod_inv.mod_mul1/_200_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_201_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_265_  (.A(\uut.mod_inv.mod_mul1/_197_ ),
    .B(\uut.mod_inv.mod_mul1/_201_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_202_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_266_  (.A(\uut.mod_inv.mod_mul1/_192_ ),
    .B(\uut.mod_inv.mod_mul1/_202_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_203_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_267_  (.A_N(\uut.sel_in_sh3.m0.Q ),
    .B(\uut.mod_inv.mod_mul1/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_204_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul1/_268_  (.A1(\uut.mod_inv.mod_mul1/_193_ ),
    .A2(\uut.mod_inv.mod_mul1/_189_ ),
    .B1_N(\uut.mod_inv.mod_mul1/_204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_205_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_269_  (.A(\uut.sel_in_sh3.m5.Q ),
    .B_N(\uut.mod_inv.mod_mul1/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_206_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_270_  (.A0(\uut.mod_inv.mod_mul1/_204_ ),
    .A1(\uut.mod_inv.mod_mul1/_205_ ),
    .S(\uut.mod_inv.mod_mul1/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_207_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_271_  (.A(\uut.mod_inv.mod_mul1/_203_ ),
    .B(\uut.mod_inv.mod_mul1/_207_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_208_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_272_  (.A(\uut.sel_in_sh1.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_209_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_273_  (.A_N(net28),
    .B(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_210_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_274_  (.A0(\uut.in1[0] ),
    .A1(net28),
    .S(\uut.sel_in_sh1.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_211_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_275_  (.A(\uut.sel_in_sh3.m6.Q ),
    .B_N(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_212_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_276_  (.A0(\uut.mod_inv.mod_mul1/_210_ ),
    .A1(\uut.mod_inv.mod_mul1/_211_ ),
    .S(\uut.mod_inv.mod_mul1/_212_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_213_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_277_  (.A_N(\uut.sel_in_sh3.m3.Q ),
    .B(\uut.sel_in_sh1.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_214_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_278_  (.A(\uut.sel_in_sh1.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_215_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_279_  (.A0(\uut.mod_inv.mod_mul1/_215_ ),
    .A1(\uut.sel_in_sh3.m3.Q ),
    .S(\uut.sel_in_sh1.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_216_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_280_  (.A(\uut.sel_in_sh3.m7.Q ),
    .B_N(\uut.sel_in_sh1.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_217_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_281_  (.A0(\uut.mod_inv.mod_mul1/_214_ ),
    .A1(\uut.mod_inv.mod_mul1/_216_ ),
    .S(\uut.mod_inv.mod_mul1/_217_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_218_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_282_  (.A(\uut.mod_inv.mod_mul1/_213_ ),
    .B(\uut.mod_inv.mod_mul1/_218_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_219_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_283_  (.A_N(\uut.sel_in_sh3.m5.Q ),
    .B(\uut.mod_inv.mod_mul1/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_220_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_284_  (.A0(\uut.sel_in_sh1.m5.Q ),
    .A1(\uut.sel_in_sh3.m5.Q ),
    .S(\uut.sel_in_sh1.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_000_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_285_  (.A(\uut.sel_in_sh3.m3.Q ),
    .B_N(\uut.sel_in_sh1.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_001_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul1/_286_  (.A0(\uut.mod_inv.mod_mul1/_220_ ),
    .A1(\uut.mod_inv.mod_mul1/_000_ ),
    .S(\uut.mod_inv.mod_mul1/_001_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_002_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_287_  (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_003_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_288_  (.A_N(\uut.sel_in_sh3.m1.Q ),
    .B(\uut.mod_inv.mod_mul1/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_004_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_289_  (.A(\uut.sel_in_sh1.m1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_005_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_290_  (.A0(\uut.mod_inv.mod_mul1/_005_ ),
    .A1(\uut.sel_in_sh3.m1.Q ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_006_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_291_  (.A(\uut.sel_in_sh3.m4.Q ),
    .B_N(\uut.mod_inv.mod_mul1/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_007_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_292_  (.A0(\uut.mod_inv.mod_mul1/_004_ ),
    .A1(\uut.mod_inv.mod_mul1/_006_ ),
    .S(\uut.mod_inv.mod_mul1/_007_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_008_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul1/_293_  (.A(\uut.mod_inv.mod_mul1/_002_ ),
    .B(\uut.mod_inv.mod_mul1/_008_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_009_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_294_  (.A(\uut.mod_inv.mod_mul1/_219_ ),
    .B(\uut.mod_inv.mod_mul1/_009_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_010_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_295_  (.A_N(\uut.sel_in_sh3.m4.Q ),
    .B(\uut.mod_inv.mod_mul1/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_011_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul1/_296_  (.A1(\uut.mod_inv.mod_mul1/_215_ ),
    .A2(\uut.mod_inv.mod_mul1/_003_ ),
    .B1_N(\uut.mod_inv.mod_mul1/_011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_012_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_297_  (.A(\uut.sel_in_sh3.m3.Q ),
    .B_N(\uut.mod_inv.mod_mul1/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_013_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_298_  (.A0(\uut.mod_inv.mod_mul1/_011_ ),
    .A1(\uut.mod_inv.mod_mul1/_012_ ),
    .S(\uut.mod_inv.mod_mul1/_013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_014_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_299_  (.A_N(\uut.sel_in_sh3.m1.Q ),
    .B(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_015_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_300_  (.A0(\uut.mod_inv.mod_mul1/_005_ ),
    .A1(\uut.sel_in_sh3.m1.Q ),
    .S(\uut.sel_in_sh1.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_016_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_301_  (.A(\uut.sel_in_sh3.m6.Q ),
    .B_N(\uut.sel_in_sh1.m1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_017_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_302_  (.A0(\uut.mod_inv.mod_mul1/_015_ ),
    .A1(\uut.mod_inv.mod_mul1/_016_ ),
    .S(\uut.mod_inv.mod_mul1/_017_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_018_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_303_  (.A_N(net28),
    .B(\uut.mod_inv.mod_mul1/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_019_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul1/_304_  (.A(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_020_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_305_  (.A0(\uut.mod_inv.mod_mul1/_020_ ),
    .A1(net28),
    .S(\uut.sel_in_sh1.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_021_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_306_  (.A(\uut.sel_in_sh3.m5.Q ),
    .B_N(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_022_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_307_  (.A0(\uut.mod_inv.mod_mul1/_019_ ),
    .A1(\uut.mod_inv.mod_mul1/_021_ ),
    .S(\uut.mod_inv.mod_mul1/_022_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_023_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_308_  (.A(\uut.mod_inv.mod_mul1/_018_ ),
    .B(\uut.mod_inv.mod_mul1/_023_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_024_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_309_  (.A(\uut.mod_inv.mod_mul1/_014_ ),
    .B(\uut.mod_inv.mod_mul1/_024_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_025_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_310_  (.A(\uut.mod_inv.mod_mul1/_010_ ),
    .B(\uut.mod_inv.mod_mul1/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_026_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_311_  (.A(\uut.mod_inv.mod_mul1/_208_ ),
    .B(\uut.mod_inv.mod_mul1/_026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out2[3] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_312_  (.A(\uut.sel_in_sh2.m1.Q ),
    .B(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_027_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_313_  (.A(\uut.sel_in_sh2.m6.Q ),
    .B(\uut.mod_inv.mod_mul1/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_028_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_314_  (.A(\uut.mod_inv.mod_mul1/_027_ ),
    .B(\uut.mod_inv.mod_mul1/_028_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_029_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_315_  (.A(\uut.sel_in_sh2.m0.Q ),
    .B(\uut.mod_inv.mod_mul1/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_030_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_316_  (.A(\uut.sel_in_sh2.m7.Q ),
    .B(\uut.mod_inv.mod_mul1/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_031_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_317_  (.A(\uut.mod_inv.mod_mul1/_030_ ),
    .B(\uut.mod_inv.mod_mul1/_031_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_032_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_318_  (.A(\uut.mod_inv.mod_mul1/_029_ ),
    .B(\uut.mod_inv.mod_mul1/_032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_033_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_319_  (.A1(\uut.sel_in_sh2.m1.Q ),
    .A2(\uut.mod_inv.mod_mul1/_187_ ),
    .B1(\uut.mod_inv.mod_mul1/_005_ ),
    .B2(\uut.sel_in_sh2.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_034_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_320_  (.A(\uut.sel_in_sh2.m7.Q ),
    .B(\uut.sel_in_sh2.m1.Q ),
    .C(\uut.mod_inv.mod_mul1/_187_ ),
    .D(\uut.mod_inv.mod_mul1/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_035_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_321_  (.A(\uut.mod_inv.mod_mul1/_034_ ),
    .B(\uut.mod_inv.mod_mul1/_035_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_036_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_322_  (.A(net27),
    .B(\uut.mod_inv.mod_mul1/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_037_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_323_  (.A(\uut.sel_in_sh2.m5.Q ),
    .B(\uut.mod_inv.mod_mul1/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_038_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_324_  (.A(\uut.mod_inv.mod_mul1/_037_ ),
    .B(\uut.mod_inv.mod_mul1/_038_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_039_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_325_  (.A(\uut.mod_inv.mod_mul1/_036_ ),
    .B(\uut.mod_inv.mod_mul1/_039_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_040_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_326_  (.A(\uut.mod_inv.mod_mul1/_033_ ),
    .B(\uut.mod_inv.mod_mul1/_040_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_041_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_327_  (.A1(\uut.sel_in_sh2.m5.Q ),
    .A2(\uut.mod_inv.mod_mul1/_215_ ),
    .B1(\uut.mod_inv.mod_mul1/_193_ ),
    .B2(\uut.sel_in_sh2.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_042_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_328_  (.A(\uut.sel_in_sh2.m3.Q ),
    .B(\uut.sel_in_sh2.m5.Q ),
    .C(\uut.mod_inv.mod_mul1/_215_ ),
    .D(\uut.mod_inv.mod_mul1/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_043_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_329_  (.A(\uut.mod_inv.mod_mul1/_042_ ),
    .B(\uut.mod_inv.mod_mul1/_043_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_044_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_330_  (.A(\uut.sel_in_sh2.m7.Q ),
    .B(\uut.mod_inv.mod_mul1/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_045_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_331_  (.A(\uut.sel_in_sh2.m3.Q ),
    .B(\uut.mod_inv.mod_mul1/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_046_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_332_  (.A(\uut.mod_inv.mod_mul1/_045_ ),
    .B(\uut.mod_inv.mod_mul1/_046_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_047_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_333_  (.A(\uut.mod_inv.mod_mul1/_044_ ),
    .B(\uut.mod_inv.mod_mul1/_047_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_048_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_334_  (.A(net12),
    .B(\uut.mod_inv.mod_mul1/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_049_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_335_  (.A(\uut.sel_in_sh2.m3.Q ),
    .B(\uut.mod_inv.mod_mul1/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_050_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_336_  (.A(\uut.mod_inv.mod_mul1/_049_ ),
    .B(\uut.mod_inv.mod_mul1/_050_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_051_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_337_  (.A(\uut.mod_inv.mod_mul1/_048_ ),
    .B(\uut.mod_inv.mod_mul1/_051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_052_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_338_  (.A1(\uut.sel_in_sh2.m1.Q ),
    .A2(\uut.mod_inv.mod_mul1/_193_ ),
    .B1(\uut.mod_inv.mod_mul1/_005_ ),
    .B2(\uut.sel_in_sh2.m5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_053_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_339_  (.A(\uut.sel_in_sh2.m5.Q ),
    .B(\uut.sel_in_sh2.m1.Q ),
    .C(\uut.mod_inv.mod_mul1/_193_ ),
    .D(\uut.mod_inv.mod_mul1/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_054_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_340_  (.A(\uut.mod_inv.mod_mul1/_053_ ),
    .B(\uut.mod_inv.mod_mul1/_054_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_055_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_341_  (.A1(\uut.sel_in_sh2.m1.Q ),
    .A2(\uut.mod_inv.mod_mul1/_003_ ),
    .B1(\uut.mod_inv.mod_mul1/_005_ ),
    .B2(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_056_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_342_  (.A(net12),
    .B(\uut.sel_in_sh2.m1.Q ),
    .C(\uut.mod_inv.mod_mul1/_003_ ),
    .D(\uut.mod_inv.mod_mul1/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_057_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_343_  (.A(\uut.mod_inv.mod_mul1/_056_ ),
    .B(\uut.mod_inv.mod_mul1/_057_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_058_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_344_  (.A(\uut.mod_inv.mod_mul1/_055_ ),
    .B(\uut.mod_inv.mod_mul1/_058_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_059_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_345_  (.A1(net27),
    .A2(\uut.mod_inv.mod_mul1/_209_ ),
    .B1(\uut.mod_inv.mod_mul1/_020_ ),
    .B2(\uut.sel_in_sh2.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_060_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_346_  (.A(\uut.sel_in_sh2.m6.Q ),
    .B(net27),
    .C(\uut.mod_inv.mod_mul1/_209_ ),
    .D(\uut.mod_inv.mod_mul1/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_061_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_347_  (.A(\uut.mod_inv.mod_mul1/_060_ ),
    .B(\uut.mod_inv.mod_mul1/_061_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_062_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_348_  (.A(\uut.sel_in_sh2.m5.Q ),
    .B(\uut.mod_inv.mod_mul1/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_063_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_349_  (.A(\uut.sel_in_sh2.m0.Q ),
    .B(\uut.mod_inv.mod_mul1/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_064_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_350_  (.A(\uut.mod_inv.mod_mul1/_063_ ),
    .B(\uut.mod_inv.mod_mul1/_064_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_065_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_351_  (.A(\uut.mod_inv.mod_mul1/_062_ ),
    .B(\uut.mod_inv.mod_mul1/_065_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_066_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_352_  (.A(\uut.mod_inv.mod_mul1/_059_ ),
    .B(\uut.mod_inv.mod_mul1/_066_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_067_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_353_  (.A(\uut.mod_inv.mod_mul1/_052_ ),
    .B(\uut.mod_inv.mod_mul1/_067_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_068_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_354_  (.A(\uut.mod_inv.mod_mul1/_041_ ),
    .B(\uut.mod_inv.mod_mul1/_068_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out3[3] ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.mod_mul1/_355_  (.A1(\uut.mod_inv.mod_mul1/_160_ ),
    .A2(\uut.mod_inv.mod_mul1/_164_ ),
    .B1_N(\uut.mod_inv.mod_mul1/_161_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_069_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_356_  (.A(\uut.mod_inv.mod_mul1/_160_ ),
    .B(\uut.mod_inv.mod_mul1/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_070_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_357_  (.A(\uut.mod_inv.mod_mul1/_162_ ),
    .B(\uut.mod_inv.mod_mul1/_070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_071_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_358_  (.A0(\uut.mod_inv.mod_mul1/_159_ ),
    .A1(\uut.mod_inv.mod_mul1/_069_ ),
    .S(\uut.mod_inv.mod_mul1/_071_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_072_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_359_  (.A(\uut.sel_in_sh3.m4.Q ),
    .B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_073_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_360_  (.A(\uut.mod_inv.mod_mul1/_163_ ),
    .B(\uut.mod_inv.mod_mul1/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_074_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul1/_361_  (.A(\uut.mod_inv.mod_mul1/_159_ ),
    .B(\uut.mod_inv.mod_mul1/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_075_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_362_  (.A(\uut.mod_inv.mod_mul1/_162_ ),
    .B(\uut.mod_inv.mod_mul1/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_076_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_363_  (.A(\uut.mod_inv.mod_mul1/_075_ ),
    .B(\uut.mod_inv.mod_mul1/_076_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_364_  (.A(\uut.mod_inv.mod_mul1/_074_ ),
    .B(\uut.mod_inv.mod_mul1/_077_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_078_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_365_  (.A(\uut.mod_inv.mod_mul1/_173_ ),
    .B(\uut.mod_inv.mod_mul1/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_079_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_366_  (.A0(\uut.mod_inv.mod_mul1/_168_ ),
    .A1(\uut.mod_inv.mod_mul1/_170_ ),
    .S(\uut.mod_inv.mod_mul1/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_080_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_367_  (.A(\uut.mod_inv.mod_mul1/_079_ ),
    .B(\uut.mod_inv.mod_mul1/_080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_081_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_368_  (.A(\uut.mod_inv.mod_mul1/_078_ ),
    .B(\uut.mod_inv.mod_mul1/_081_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_082_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_369_  (.A(\uut.mod_inv.mod_mul1/_072_ ),
    .B(\uut.mod_inv.mod_mul1/_082_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out1[2] ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_370_  (.A_N(net28),
    .B(\uut.mod_inv.mod_mul1/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_083_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_371_  (.A0(\uut.mod_inv.mod_mul1/_020_ ),
    .A1(net28),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_084_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_372_  (.A(\uut.sel_in_sh3.m4.Q ),
    .B_N(\uut.in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_085_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_373_  (.A0(\uut.mod_inv.mod_mul1/_083_ ),
    .A1(\uut.mod_inv.mod_mul1/_084_ ),
    .S(\uut.mod_inv.mod_mul1/_085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_086_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_374_  (.A(\uut.mod_inv.mod_mul1/_201_ ),
    .B(\uut.mod_inv.mod_mul1/_086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_087_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_375_  (.A_N(\uut.sel_in_sh3.m0.Q ),
    .B(\uut.sel_in_sh1.m4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_088_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_376_  (.A0(\uut.sel_in_sh1.m0.Q ),
    .A1(\uut.sel_in_sh3.m0.Q ),
    .S(\uut.sel_in_sh1.m4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_089_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_377_  (.A(\uut.sel_in_sh3.m4.Q ),
    .B_N(\uut.sel_in_sh1.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_090_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_378_  (.A0(\uut.mod_inv.mod_mul1/_088_ ),
    .A1(\uut.mod_inv.mod_mul1/_089_ ),
    .S(\uut.mod_inv.mod_mul1/_090_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_091_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_379_  (.A_N(\uut.sel_in_sh3.m0.Q ),
    .B(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_092_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_380_  (.A0(\uut.mod_inv.mod_mul1/_189_ ),
    .A1(\uut.sel_in_sh3.m0.Q ),
    .S(\uut.sel_in_sh1.m6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_093_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_381_  (.A(\uut.sel_in_sh3.m6.Q ),
    .B_N(\uut.sel_in_sh1.m0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_094_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_382_  (.A0(\uut.mod_inv.mod_mul1/_092_ ),
    .A1(\uut.mod_inv.mod_mul1/_093_ ),
    .S(\uut.mod_inv.mod_mul1/_094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_095_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_383_  (.A(\uut.mod_inv.mod_mul1/_091_ ),
    .B(\uut.mod_inv.mod_mul1/_095_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_096_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_384_  (.A(\uut.mod_inv.mod_mul1/_087_ ),
    .B(\uut.mod_inv.mod_mul1/_096_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_097_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_385_  (.A_N(net28),
    .B(\uut.mod_inv.mod_mul1/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_098_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul1/_386_  (.A1(\uut.mod_inv.mod_mul1/_187_ ),
    .A2(\uut.mod_inv.mod_mul1/_020_ ),
    .B1_N(\uut.mod_inv.mod_mul1/_098_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_099_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_387_  (.A(\uut.sel_in_sh3.m7.Q ),
    .B_N(\uut.mod_inv.mod_mul1/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_100_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_388_  (.A0(\uut.mod_inv.mod_mul1/_098_ ),
    .A1(\uut.mod_inv.mod_mul1/_099_ ),
    .S(\uut.mod_inv.mod_mul1/_100_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_101_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul1/_389_  (.A_N(\uut.sel_in_sh3.m6.Q ),
    .B(\uut.mod_inv.mod_mul1/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_102_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_390_  (.A0(\uut.mod_inv.mod_mul1/_209_ ),
    .A1(\uut.sel_in_sh3.m6.Q ),
    .S(\uut.sel_in_sh1.m3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_103_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul1/_391_  (.A(\uut.sel_in_sh3.m3.Q ),
    .B_N(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_104_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_392_  (.A0(\uut.mod_inv.mod_mul1/_102_ ),
    .A1(\uut.mod_inv.mod_mul1/_103_ ),
    .S(\uut.mod_inv.mod_mul1/_104_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_105_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_393_  (.A(\uut.mod_inv.mod_mul1/_002_ ),
    .B(\uut.mod_inv.mod_mul1/_105_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_106_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_394_  (.A(\uut.mod_inv.mod_mul1/_101_ ),
    .B(\uut.mod_inv.mod_mul1/_106_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_107_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_395_  (.A(\uut.mod_inv.mod_mul1/_197_ ),
    .B(\uut.mod_inv.mod_mul1/_213_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_108_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_396_  (.A(\uut.mod_inv.mod_mul1/_107_ ),
    .B(\uut.mod_inv.mod_mul1/_108_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_109_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_397_  (.A(\uut.mod_inv.mod_mul1/_097_ ),
    .B(\uut.mod_inv.mod_mul1/_109_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out2[2] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_398_  (.A(\uut.sel_in_sh2.m6.Q ),
    .B(\uut.mod_inv.mod_mul1/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_110_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_399_  (.A(\uut.mod_inv.mod_mul1/_055_ ),
    .B(\uut.mod_inv.mod_mul1/_110_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_111_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_400_  (.A(\uut.sel_in_sh2.m3.Q ),
    .B(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_112_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_401_  (.A1(net27),
    .A2(\uut.mod_inv.mod_mul1/_187_ ),
    .B1(\uut.mod_inv.mod_mul1/_020_ ),
    .B2(\uut.sel_in_sh2.m7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_113_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_402_  (.A(\uut.sel_in_sh2.m7.Q ),
    .B(net27),
    .C(\uut.mod_inv.mod_mul1/_187_ ),
    .D(\uut.mod_inv.mod_mul1/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_114_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_403_  (.A(\uut.mod_inv.mod_mul1/_113_ ),
    .B(\uut.mod_inv.mod_mul1/_114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_115_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_404_  (.A(\uut.mod_inv.mod_mul1/_112_ ),
    .B(\uut.mod_inv.mod_mul1/_115_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_116_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_405_  (.A(\uut.mod_inv.mod_mul1/_111_ ),
    .B(\uut.mod_inv.mod_mul1/_116_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_117_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_406_  (.A(\uut.mod_inv.mod_mul1/_044_ ),
    .B(\uut.mod_inv.mod_mul1/_117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_118_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_407_  (.A(\uut.sel_in_sh2.m6.Q ),
    .B(\uut.mod_inv.mod_mul1/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_119_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_408_  (.A(\uut.sel_in_sh2.m0.Q ),
    .B(\uut.mod_inv.mod_mul1/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_120_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_409_  (.A(\uut.mod_inv.mod_mul1/_119_ ),
    .B(\uut.mod_inv.mod_mul1/_120_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_121_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_410_  (.A(\uut.mod_inv.mod_mul1/_036_ ),
    .B(\uut.mod_inv.mod_mul1/_121_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_122_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_411_  (.A(\uut.mod_inv.mod_mul1/_062_ ),
    .B(\uut.mod_inv.mod_mul1/_122_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_123_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul1/_412_  (.A1(\uut.sel_in_sh2.m0.Q ),
    .A2(\uut.mod_inv.mod_mul1/_003_ ),
    .B1(\uut.mod_inv.mod_mul1/_189_ ),
    .B2(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_124_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul1/_413_  (.A(net12),
    .B(\uut.sel_in_sh2.m0.Q ),
    .C(\uut.mod_inv.mod_mul1/_003_ ),
    .D(\uut.mod_inv.mod_mul1/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_125_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_414_  (.A(\uut.mod_inv.mod_mul1/_124_ ),
    .B(\uut.mod_inv.mod_mul1/_125_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_126_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_415_  (.A(\uut.sel_in_sh2.m4.Q ),
    .B(\uut.mod_inv.mod_mul1/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_127_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_416_  (.A(net27),
    .B(\uut.mod_inv.mod_mul1/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_128_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_417_  (.A(\uut.mod_inv.mod_mul1/_127_ ),
    .B(\uut.mod_inv.mod_mul1/_128_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_129_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_418_  (.A(\uut.mod_inv.mod_mul1/_126_ ),
    .B(\uut.mod_inv.mod_mul1/_129_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_130_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_419_  (.A(\uut.mod_inv.mod_mul1/_123_ ),
    .B(\uut.mod_inv.mod_mul1/_130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_131_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_420_  (.A(\uut.mod_inv.mod_mul1/_118_ ),
    .B(\uut.mod_inv.mod_mul1/_131_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out3[2] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_421_  (.A(\uut.mod_inv.mod_mul1/_075_ ),
    .B(\uut.mod_inv.mod_mul1/_079_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_132_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul1/_422_  (.A(\uut.mod_inv.mod_mul1/_163_ ),
    .B(\uut.mod_inv.mod_mul1/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_133_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.mod_mul1/_423_  (.A(\uut.mod_inv.mod_mul1/_166_ ),
    .B(\uut.mod_inv.mod_mul1/_169_ ),
    .C(\uut.mod_inv.mod_mul1/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_134_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.mod_mul1/_424_  (.A(\uut.mod_inv.mod_mul1/_166_ ),
    .B(\uut.mod_inv.mod_mul1/_167_ ),
    .C(\uut.mod_inv.mod_mul1/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_135_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_425_  (.A(\uut.mod_inv.mod_mul1/_163_ ),
    .B(\uut.mod_inv.mod_mul1/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_136_ ));
 sky130_fd_sc_hd__a32o_1 \uut.mod_inv.mod_mul1/_426_  (.A1(\uut.mod_inv.mod_mul1/_133_ ),
    .A2(\uut.mod_inv.mod_mul1/_134_ ),
    .A3(\uut.mod_inv.mod_mul1/_135_ ),
    .B1(\uut.mod_inv.mod_mul1/_136_ ),
    .B2(\uut.mod_inv.mod_mul1/_170_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_137_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_427_  (.A(\uut.mod_inv.mod_mul1/_179_ ),
    .B(\uut.mod_inv.mod_mul1/_137_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_138_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.mod_mul1/_428_  (.A(\uut.mod_inv.mod_mul1/_162_ ),
    .B(\uut.mod_inv.mod_mul1/_166_ ),
    .C_N(\uut.mod_inv.mod_mul1/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_139_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul1/_429_  (.A(\uut.mod_inv.mod_mul1/_161_ ),
    .B(\uut.mod_inv.mod_mul1/_139_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_140_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.mod_mul1/_430_  (.A(\uut.mod_inv.mod_mul1/_160_ ),
    .B(\uut.mod_inv.mod_mul1/_166_ ),
    .C_N(\uut.mod_inv.mod_mul1/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_141_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_431_  (.A0(\uut.mod_inv.mod_mul1/_163_ ),
    .A1(\uut.mod_inv.mod_mul1/_070_ ),
    .S(\uut.mod_inv.mod_mul1/_141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_142_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul1/_432_  (.A0(\uut.mod_inv.mod_mul1/_140_ ),
    .A1(\uut.mod_inv.mod_mul1/_161_ ),
    .S(\uut.mod_inv.mod_mul1/_142_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_143_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_433_  (.A(\uut.mod_inv.mod_mul1/_138_ ),
    .B(\uut.mod_inv.mod_mul1/_143_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_144_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_434_  (.A(\uut.mod_inv.mod_mul1/_132_ ),
    .B(\uut.mod_inv.mod_mul1/_144_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out1[1] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_435_  (.A(\uut.mod_inv.mod_mul1/_203_ ),
    .B(\uut.mod_inv.mod_mul1/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_145_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_436_  (.A(\uut.mod_inv.mod_mul1/_218_ ),
    .B(\uut.mod_inv.mod_mul1/_091_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_146_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_437_  (.A(\uut.mod_inv.mod_mul1/_107_ ),
    .B(\uut.mod_inv.mod_mul1/_146_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_147_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_438_  (.A(\uut.mod_inv.mod_mul1/_145_ ),
    .B(\uut.mod_inv.mod_mul1/_147_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out2[1] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_439_  (.A(\uut.mod_inv.mod_mul1/_052_ ),
    .B(\uut.mod_inv.mod_mul1/_126_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_148_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_440_  (.A(\uut.mod_inv.mod_mul1/_041_ ),
    .B(\uut.mod_inv.mod_mul1/_117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_149_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_441_  (.A(\uut.mod_inv.mod_mul1/_148_ ),
    .B(\uut.mod_inv.mod_mul1/_149_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out3[1] ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.mod_mul1/_442_  (.A1(\uut.mod_inv.mod_mul1/_162_ ),
    .A2(\uut.mod_inv.mod_mul1/_079_ ),
    .B1(\uut.mod_inv.mod_mul1/_076_ ),
    .B2(\uut.mod_inv.mod_mul1/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_150_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul1/_443_  (.A(\uut.mod_inv.mod_mul1/_159_ ),
    .B(\uut.mod_inv.mod_mul1/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_151_ ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.mod_mul1/_444_  (.A1(\uut.mod_inv.mod_mul1/_163_ ),
    .A2(\uut.mod_inv.mod_mul1/_151_ ),
    .B1(\uut.mod_inv.mod_mul1/_074_ ),
    .B2(\uut.mod_inv.mod_mul1/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_152_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_445_  (.A(\uut.mod_inv.mod_mul1/_150_ ),
    .B(\uut.mod_inv.mod_mul1/_152_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_153_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_446_  (.A(\uut.mod_inv.mod_mul1/_175_ ),
    .B(\uut.mod_inv.mod_mul1/_153_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_154_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_447_  (.A(\uut.mod_inv.mod_mul1/_172_ ),
    .B(\uut.mod_inv.mod_mul1/_154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out1[0] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul1/_448_  (.A(\uut.mod_inv.mod_mul1/_207_ ),
    .B(\uut.mod_inv.mod_mul1/_097_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul1/_155_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_449_  (.A(\uut.mod_inv.mod_mul1/_010_ ),
    .B(\uut.mod_inv.mod_mul1/_155_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out2[0] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_450_  (.A(\uut.mod_inv.mod_mul1/_058_ ),
    .B(\uut.mod_inv.mod_mul1/_130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_156_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul1/_451_  (.A(\uut.mod_inv.mod_mul1/_066_ ),
    .B(\uut.mod_inv.mod_mul1/_122_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_157_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_452_  (.A(\uut.mod_inv.mod_mul1/_156_ ),
    .B(\uut.mod_inv.mod_mul1/_157_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1/_158_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul1/_453_  (.A(\uut.mod_inv.mod_mul1/_048_ ),
    .B(\uut.mod_inv.mod_mul1/_158_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul1_out3[0] ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_221_  (.A(net17),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_159_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_222_  (.A(\uut.mod_inv.sh3_reg_1_1[3] ),
    .B(\uut.mod_inv.sh2_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_160_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul2/_223_  (.A(\uut.mod_inv.mod_mul2/_159_ ),
    .B(\uut.mod_inv.mod_mul2/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_161_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_224_  (.A(\uut.mod_inv.sh3_reg_1_1[2] ),
    .B(\uut.mod_inv.sh2_reg_1_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_162_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_225_  (.A(net15),
    .B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_163_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_226_  (.A(\uut.mod_inv.mod_mul2/_162_ ),
    .B(\uut.mod_inv.mod_mul2/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_164_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_227_  (.A(\uut.mod_inv.mod_mul2/_161_ ),
    .B(\uut.mod_inv.mod_mul2/_164_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_165_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_228_  (.A(net14),
    .B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_166_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul2/_229_  (.A(\uut.mod_inv.sh3_reg_1_1[1] ),
    .B(\uut.mod_inv.sh2_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_167_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_230_  (.A(\uut.mod_inv.mod_mul2/_166_ ),
    .B(\uut.mod_inv.mod_mul2/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_168_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_231_  (.A(\uut.mod_inv.sh3_reg_1_1[1] ),
    .B(\uut.mod_inv.sh2_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_169_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_232_  (.A(\uut.mod_inv.mod_mul2/_166_ ),
    .B(\uut.mod_inv.mod_mul2/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_170_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_233_  (.A0(\uut.mod_inv.mod_mul2/_168_ ),
    .A1(\uut.mod_inv.mod_mul2/_170_ ),
    .S(\uut.mod_inv.mod_mul2/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_171_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_234_  (.A(\uut.mod_inv.mod_mul2/_165_ ),
    .B(\uut.mod_inv.mod_mul2/_171_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_172_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_235_  (.A(net19),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_173_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_236_  (.A(\uut.mod_inv.mod_mul2/_167_ ),
    .B(\uut.mod_inv.mod_mul2/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_174_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul2/_237_  (.A(\uut.mod_inv.mod_mul2/_169_ ),
    .B(\uut.mod_inv.mod_mul2/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_175_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_238_  (.A0(\uut.mod_inv.mod_mul2/_174_ ),
    .A1(\uut.mod_inv.mod_mul2/_175_ ),
    .S(\uut.mod_inv.mod_mul2/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_176_ ));
 sky130_fd_sc_hd__o22a_1 \uut.mod_inv.mod_mul2/_239_  (.A1(\uut.mod_inv.mod_mul2/_159_ ),
    .A2(\uut.mod_inv.mod_mul2/_162_ ),
    .B1(\uut.mod_inv.mod_mul2/_173_ ),
    .B2(\uut.mod_inv.mod_mul2/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_177_ ));
 sky130_fd_sc_hd__or4_1 \uut.mod_inv.mod_mul2/_240_  (.A(\uut.mod_inv.mod_mul2/_159_ ),
    .B(\uut.mod_inv.mod_mul2/_160_ ),
    .C(\uut.mod_inv.mod_mul2/_162_ ),
    .D(\uut.mod_inv.mod_mul2/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_178_ ));
 sky130_fd_sc_hd__nor2b_1 \uut.mod_inv.mod_mul2/_241_  (.A(\uut.mod_inv.mod_mul2/_177_ ),
    .B_N(\uut.mod_inv.mod_mul2/_178_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_179_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_242_  (.A(\uut.mod_inv.mod_mul2/_159_ ),
    .B(\uut.mod_inv.mod_mul2/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_180_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_243_  (.A(\uut.mod_inv.sh3_reg_1_1[0] ),
    .B(\uut.mod_inv.sh2_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_181_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_244_  (.A0(\uut.mod_inv.mod_mul2/_167_ ),
    .A1(\uut.mod_inv.mod_mul2/_181_ ),
    .S(\uut.mod_inv.mod_mul2/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_182_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_245_  (.A(\uut.mod_inv.mod_mul2/_166_ ),
    .B(\uut.mod_inv.mod_mul2/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_183_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_246_  (.A0(\uut.mod_inv.mod_mul2/_180_ ),
    .A1(\uut.mod_inv.mod_mul2/_182_ ),
    .S(\uut.mod_inv.mod_mul2/_183_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_184_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_247_  (.A(\uut.mod_inv.mod_mul2/_179_ ),
    .B(\uut.mod_inv.mod_mul2/_184_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_185_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_248_  (.A(\uut.mod_inv.mod_mul2/_176_ ),
    .B(\uut.mod_inv.mod_mul2/_185_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_186_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_249_  (.A(\uut.mod_inv.mod_mul2/_172_ ),
    .B(\uut.mod_inv.mod_mul2/_186_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out1[3] ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_250_  (.A(\uut.mod_inv.sh1_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_187_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_251_  (.A_N(net19),
    .B(\uut.mod_inv.mod_mul2/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_188_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_252_  (.A(\uut.mod_inv.mul_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_189_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul2/_253_  (.A1(\uut.mod_inv.mod_mul2/_187_ ),
    .A2(\uut.mod_inv.mod_mul2/_189_ ),
    .B1_N(\uut.mod_inv.mod_mul2/_188_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_190_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_254_  (.A(\uut.mod_inv.sh3_reg_1_1[3] ),
    .B_N(\uut.mod_inv.mod_mul2/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_191_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_255_  (.A0(\uut.mod_inv.mod_mul2/_188_ ),
    .A1(\uut.mod_inv.mod_mul2/_190_ ),
    .S(\uut.mod_inv.mod_mul2/_191_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_192_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_256_  (.A(\uut.mod_inv.sh1_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_193_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_257_  (.A_N(net17),
    .B(\uut.mod_inv.mod_mul2/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_194_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_258_  (.A0(net20),
    .A1(net17),
    .S(\uut.mod_inv.sh1_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_195_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_259_  (.A(\uut.mod_inv.sh3_reg_1_1[1] ),
    .B_N(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_196_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_260_  (.A0(\uut.mod_inv.mod_mul2/_194_ ),
    .A1(\uut.mod_inv.mod_mul2/_195_ ),
    .S(\uut.mod_inv.mod_mul2/_196_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_197_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_261_  (.A_N(net17),
    .B(\uut.mod_inv.sh1_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_198_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_262_  (.A0(net20),
    .A1(net17),
    .S(\uut.mod_inv.sh1_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_199_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_263_  (.A(\uut.mod_inv.sh3_reg_1_1[3] ),
    .B_N(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_200_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_264_  (.A0(\uut.mod_inv.mod_mul2/_198_ ),
    .A1(\uut.mod_inv.mod_mul2/_199_ ),
    .S(\uut.mod_inv.mod_mul2/_200_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_201_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_265_  (.A(\uut.mod_inv.mod_mul2/_197_ ),
    .B(\uut.mod_inv.mod_mul2/_201_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_202_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_266_  (.A(\uut.mod_inv.mod_mul2/_192_ ),
    .B(\uut.mod_inv.mod_mul2/_202_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_203_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_267_  (.A_N(net19),
    .B(\uut.mod_inv.mod_mul2/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_204_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul2/_268_  (.A1(\uut.mod_inv.mod_mul2/_193_ ),
    .A2(\uut.mod_inv.mod_mul2/_189_ ),
    .B1_N(\uut.mod_inv.mod_mul2/_204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_205_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_269_  (.A(\uut.mod_inv.sh3_reg_1_1[1] ),
    .B_N(\uut.mod_inv.mod_mul2/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_206_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_270_  (.A0(\uut.mod_inv.mod_mul2/_204_ ),
    .A1(\uut.mod_inv.mod_mul2/_205_ ),
    .S(\uut.mod_inv.mod_mul2/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_207_ ));
 sky130_fd_sc_hd__xor2_4 \uut.mod_inv.mod_mul2/_271_  (.A(\uut.mod_inv.mod_mul2/_203_ ),
    .B(\uut.mod_inv.mod_mul2/_207_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_208_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_272_  (.A(\uut.mod_inv.sh1_reg_1_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_209_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_273_  (.A_N(net15),
    .B(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_210_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_274_  (.A0(\uut.mod_inv.mul_in1[2] ),
    .A1(net15),
    .S(\uut.mod_inv.sh1_reg_1_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_211_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_275_  (.A(\uut.mod_inv.sh3_reg_1_1[2] ),
    .B_N(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_212_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_276_  (.A0(\uut.mod_inv.mod_mul2/_210_ ),
    .A1(\uut.mod_inv.mod_mul2/_211_ ),
    .S(\uut.mod_inv.mod_mul2/_212_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_213_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_277_  (.A_N(net14),
    .B(\uut.mod_inv.sh1_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_214_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_278_  (.A(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_215_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_279_  (.A0(\uut.mod_inv.mod_mul2/_215_ ),
    .A1(net14),
    .S(\uut.mod_inv.sh1_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_216_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_280_  (.A(\uut.mod_inv.sh3_reg_1_1[3] ),
    .B_N(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_217_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_281_  (.A0(\uut.mod_inv.mod_mul2/_214_ ),
    .A1(\uut.mod_inv.mod_mul2/_216_ ),
    .S(\uut.mod_inv.mod_mul2/_217_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_218_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_282_  (.A(\uut.mod_inv.mod_mul2/_213_ ),
    .B(\uut.mod_inv.mod_mul2/_218_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_219_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_283_  (.A_N(\uut.mod_inv.sh3_reg_1_1[1] ),
    .B(\uut.mod_inv.mod_mul2/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_220_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_284_  (.A0(\uut.mod_inv.sh1_reg_1_1[1] ),
    .A1(\uut.mod_inv.sh3_reg_1_1[1] ),
    .S(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_000_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_285_  (.A(net14),
    .B_N(\uut.mod_inv.sh1_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_001_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_286_  (.A0(\uut.mod_inv.mod_mul2/_220_ ),
    .A1(\uut.mod_inv.mod_mul2/_000_ ),
    .S(\uut.mod_inv.mod_mul2/_001_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_002_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_287_  (.A(\uut.mod_inv.sh1_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_003_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_288_  (.A_N(net17),
    .B(\uut.mod_inv.mod_mul2/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_004_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_289_  (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_005_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_290_  (.A0(\uut.mod_inv.mod_mul2/_005_ ),
    .A1(net17),
    .S(\uut.mod_inv.sh1_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_006_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_291_  (.A(\uut.mod_inv.sh3_reg_1_1[0] ),
    .B_N(\uut.mod_inv.mod_mul2/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_007_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_292_  (.A0(\uut.mod_inv.mod_mul2/_004_ ),
    .A1(\uut.mod_inv.mod_mul2/_006_ ),
    .S(\uut.mod_inv.mod_mul2/_007_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_008_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul2/_293_  (.A(\uut.mod_inv.mod_mul2/_002_ ),
    .B(\uut.mod_inv.mod_mul2/_008_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_009_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_294_  (.A(\uut.mod_inv.mod_mul2/_219_ ),
    .B(\uut.mod_inv.mod_mul2/_009_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_010_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_295_  (.A_N(\uut.mod_inv.sh3_reg_1_1[0] ),
    .B(\uut.mod_inv.mod_mul2/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_011_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul2/_296_  (.A1(\uut.mod_inv.mod_mul2/_215_ ),
    .A2(\uut.mod_inv.mod_mul2/_003_ ),
    .B1_N(\uut.mod_inv.mod_mul2/_011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_012_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_297_  (.A(net14),
    .B_N(\uut.mod_inv.mod_mul2/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_013_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul2/_298_  (.A0(\uut.mod_inv.mod_mul2/_011_ ),
    .A1(\uut.mod_inv.mod_mul2/_012_ ),
    .S(\uut.mod_inv.mod_mul2/_013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_014_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_299_  (.A_N(net17),
    .B(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_015_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_300_  (.A0(\uut.mod_inv.mod_mul2/_005_ ),
    .A1(net17),
    .S(\uut.mod_inv.sh1_reg_1_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_016_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_301_  (.A(\uut.mod_inv.sh3_reg_1_1[2] ),
    .B_N(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_017_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_302_  (.A0(\uut.mod_inv.mod_mul2/_015_ ),
    .A1(\uut.mod_inv.mod_mul2/_016_ ),
    .S(\uut.mod_inv.mod_mul2/_017_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_018_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_303_  (.A_N(net15),
    .B(\uut.mod_inv.mod_mul2/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_019_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul2/_304_  (.A(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_020_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_305_  (.A0(\uut.mod_inv.mod_mul2/_020_ ),
    .A1(net15),
    .S(\uut.mod_inv.sh1_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_021_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_306_  (.A(\uut.mod_inv.sh3_reg_1_1[1] ),
    .B_N(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_022_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_307_  (.A0(\uut.mod_inv.mod_mul2/_019_ ),
    .A1(\uut.mod_inv.mod_mul2/_021_ ),
    .S(\uut.mod_inv.mod_mul2/_022_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_023_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_308_  (.A(\uut.mod_inv.mod_mul2/_018_ ),
    .B(\uut.mod_inv.mod_mul2/_023_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_024_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_309_  (.A(\uut.mod_inv.mod_mul2/_014_ ),
    .B(\uut.mod_inv.mod_mul2/_024_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_025_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_310_  (.A(\uut.mod_inv.mod_mul2/_010_ ),
    .B(\uut.mod_inv.mod_mul2/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_026_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_311_  (.A(\uut.mod_inv.mod_mul2/_208_ ),
    .B(\uut.mod_inv.mod_mul2/_026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out2[3] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_312_  (.A(net24),
    .B(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_027_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_313_  (.A(\uut.mod_inv.sh2_reg_1_1[2] ),
    .B(\uut.mod_inv.mod_mul2/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_028_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_314_  (.A(\uut.mod_inv.mod_mul2/_027_ ),
    .B(\uut.mod_inv.mod_mul2/_028_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_029_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_315_  (.A(net26),
    .B(\uut.mod_inv.mod_mul2/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_030_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_316_  (.A(\uut.mod_inv.sh2_reg_1_1[3] ),
    .B(\uut.mod_inv.mod_mul2/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_031_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_317_  (.A(\uut.mod_inv.mod_mul2/_030_ ),
    .B(\uut.mod_inv.mod_mul2/_031_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_032_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_318_  (.A(\uut.mod_inv.mod_mul2/_029_ ),
    .B(\uut.mod_inv.mod_mul2/_032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_033_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_319_  (.A1(net24),
    .A2(\uut.mod_inv.mod_mul2/_187_ ),
    .B1(\uut.mod_inv.mod_mul2/_005_ ),
    .B2(\uut.mod_inv.sh2_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_034_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_320_  (.A(\uut.mod_inv.sh2_reg_1_1[3] ),
    .B(net24),
    .C(\uut.mod_inv.mod_mul2/_187_ ),
    .D(\uut.mod_inv.mod_mul2/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_035_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_321_  (.A(\uut.mod_inv.mod_mul2/_034_ ),
    .B(\uut.mod_inv.mod_mul2/_035_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_036_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_322_  (.A(net23),
    .B(\uut.mod_inv.mod_mul2/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_037_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_323_  (.A(\uut.mod_inv.sh2_reg_1_1[1] ),
    .B(\uut.mod_inv.mod_mul2/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_038_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_324_  (.A(\uut.mod_inv.mod_mul2/_037_ ),
    .B(\uut.mod_inv.mod_mul2/_038_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_039_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_325_  (.A(\uut.mod_inv.mod_mul2/_036_ ),
    .B(\uut.mod_inv.mod_mul2/_039_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_040_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_326_  (.A(\uut.mod_inv.mod_mul2/_033_ ),
    .B(\uut.mod_inv.mod_mul2/_040_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_041_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_327_  (.A1(\uut.mod_inv.sh2_reg_1_1[1] ),
    .A2(\uut.mod_inv.mod_mul2/_215_ ),
    .B1(\uut.mod_inv.mod_mul2/_193_ ),
    .B2(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_042_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_328_  (.A(net22),
    .B(\uut.mod_inv.sh2_reg_1_1[1] ),
    .C(\uut.mod_inv.mod_mul2/_215_ ),
    .D(\uut.mod_inv.mod_mul2/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_043_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_329_  (.A(\uut.mod_inv.mod_mul2/_042_ ),
    .B(\uut.mod_inv.mod_mul2/_043_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_044_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_330_  (.A(\uut.mod_inv.sh2_reg_1_1[3] ),
    .B(\uut.mod_inv.mod_mul2/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_045_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_331_  (.A(net22),
    .B(\uut.mod_inv.mod_mul2/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_046_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_332_  (.A(\uut.mod_inv.mod_mul2/_045_ ),
    .B(\uut.mod_inv.mod_mul2/_046_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_047_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_333_  (.A(\uut.mod_inv.mod_mul2/_044_ ),
    .B(\uut.mod_inv.mod_mul2/_047_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_048_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_334_  (.A(\uut.mod_inv.sh2_reg_1_1[0] ),
    .B(\uut.mod_inv.mod_mul2/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_049_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_335_  (.A(net22),
    .B(\uut.mod_inv.mod_mul2/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_050_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_336_  (.A(\uut.mod_inv.mod_mul2/_049_ ),
    .B(\uut.mod_inv.mod_mul2/_050_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_051_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_337_  (.A(\uut.mod_inv.mod_mul2/_048_ ),
    .B(\uut.mod_inv.mod_mul2/_051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_052_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_338_  (.A1(net24),
    .A2(\uut.mod_inv.mod_mul2/_193_ ),
    .B1(\uut.mod_inv.mod_mul2/_005_ ),
    .B2(\uut.mod_inv.sh2_reg_1_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_053_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_339_  (.A(\uut.mod_inv.sh2_reg_1_1[1] ),
    .B(net24),
    .C(\uut.mod_inv.mod_mul2/_193_ ),
    .D(\uut.mod_inv.mod_mul2/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_054_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_340_  (.A(\uut.mod_inv.mod_mul2/_053_ ),
    .B(\uut.mod_inv.mod_mul2/_054_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_055_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_341_  (.A1(net24),
    .A2(\uut.mod_inv.mod_mul2/_003_ ),
    .B1(\uut.mod_inv.mod_mul2/_005_ ),
    .B2(\uut.mod_inv.sh2_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_056_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_342_  (.A(\uut.mod_inv.sh2_reg_1_1[0] ),
    .B(net24),
    .C(\uut.mod_inv.mod_mul2/_003_ ),
    .D(\uut.mod_inv.mod_mul2/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_057_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_343_  (.A(\uut.mod_inv.mod_mul2/_056_ ),
    .B(\uut.mod_inv.mod_mul2/_057_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_058_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_344_  (.A(\uut.mod_inv.mod_mul2/_055_ ),
    .B(\uut.mod_inv.mod_mul2/_058_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_059_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_345_  (.A1(net23),
    .A2(\uut.mod_inv.mod_mul2/_209_ ),
    .B1(\uut.mod_inv.mod_mul2/_020_ ),
    .B2(\uut.mod_inv.sh2_reg_1_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_060_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_346_  (.A(\uut.mod_inv.sh2_reg_1_1[2] ),
    .B(net23),
    .C(\uut.mod_inv.mod_mul2/_209_ ),
    .D(\uut.mod_inv.mod_mul2/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_061_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_347_  (.A(\uut.mod_inv.mod_mul2/_060_ ),
    .B(\uut.mod_inv.mod_mul2/_061_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_062_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_348_  (.A(\uut.mod_inv.sh2_reg_1_1[1] ),
    .B(\uut.mod_inv.mod_mul2/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_063_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_349_  (.A(net26),
    .B(\uut.mod_inv.mod_mul2/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_064_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_350_  (.A(\uut.mod_inv.mod_mul2/_063_ ),
    .B(\uut.mod_inv.mod_mul2/_064_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_065_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_351_  (.A(\uut.mod_inv.mod_mul2/_062_ ),
    .B(\uut.mod_inv.mod_mul2/_065_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_066_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_352_  (.A(\uut.mod_inv.mod_mul2/_059_ ),
    .B(\uut.mod_inv.mod_mul2/_066_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_067_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_353_  (.A(\uut.mod_inv.mod_mul2/_052_ ),
    .B(\uut.mod_inv.mod_mul2/_067_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_068_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_354_  (.A(\uut.mod_inv.mod_mul2/_041_ ),
    .B(\uut.mod_inv.mod_mul2/_068_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out3[3] ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.mod_mul2/_355_  (.A1(\uut.mod_inv.mod_mul2/_160_ ),
    .A2(\uut.mod_inv.mod_mul2/_164_ ),
    .B1_N(\uut.mod_inv.mod_mul2/_161_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_069_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_356_  (.A(\uut.mod_inv.mod_mul2/_160_ ),
    .B(\uut.mod_inv.mod_mul2/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_070_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_357_  (.A(\uut.mod_inv.mod_mul2/_162_ ),
    .B(\uut.mod_inv.mod_mul2/_070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_071_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_358_  (.A0(\uut.mod_inv.mod_mul2/_159_ ),
    .A1(\uut.mod_inv.mod_mul2/_069_ ),
    .S(\uut.mod_inv.mod_mul2/_071_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_072_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_359_  (.A(\uut.mod_inv.sh3_reg_1_1[0] ),
    .B(\uut.mod_inv.sh2_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_073_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_360_  (.A(\uut.mod_inv.mod_mul2/_163_ ),
    .B(\uut.mod_inv.mod_mul2/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_074_ ));
 sky130_fd_sc_hd__or2_2 \uut.mod_inv.mod_mul2/_361_  (.A(\uut.mod_inv.mod_mul2/_159_ ),
    .B(\uut.mod_inv.mod_mul2/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_075_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_362_  (.A(\uut.mod_inv.mod_mul2/_162_ ),
    .B(\uut.mod_inv.mod_mul2/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_076_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_363_  (.A(\uut.mod_inv.mod_mul2/_075_ ),
    .B(\uut.mod_inv.mod_mul2/_076_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_364_  (.A(\uut.mod_inv.mod_mul2/_074_ ),
    .B(\uut.mod_inv.mod_mul2/_077_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_078_ ));
 sky130_fd_sc_hd__nor2_2 \uut.mod_inv.mod_mul2/_365_  (.A(\uut.mod_inv.mod_mul2/_173_ ),
    .B(\uut.mod_inv.mod_mul2/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_079_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_366_  (.A0(\uut.mod_inv.mod_mul2/_168_ ),
    .A1(\uut.mod_inv.mod_mul2/_170_ ),
    .S(\uut.mod_inv.mod_mul2/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_080_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_367_  (.A(\uut.mod_inv.mod_mul2/_079_ ),
    .B(\uut.mod_inv.mod_mul2/_080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_081_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_368_  (.A(\uut.mod_inv.mod_mul2/_078_ ),
    .B(\uut.mod_inv.mod_mul2/_081_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_082_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_369_  (.A(\uut.mod_inv.mod_mul2/_072_ ),
    .B(\uut.mod_inv.mod_mul2/_082_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out1[2] ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_370_  (.A_N(net15),
    .B(\uut.mod_inv.mod_mul2/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_083_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_371_  (.A0(\uut.mod_inv.mod_mul2/_020_ ),
    .A1(net15),
    .S(\uut.mod_inv.sh1_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_084_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_372_  (.A(\uut.mod_inv.sh3_reg_1_1[0] ),
    .B_N(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_085_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_373_  (.A0(\uut.mod_inv.mod_mul2/_083_ ),
    .A1(\uut.mod_inv.mod_mul2/_084_ ),
    .S(\uut.mod_inv.mod_mul2/_085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_086_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_374_  (.A(\uut.mod_inv.mod_mul2/_201_ ),
    .B(\uut.mod_inv.mod_mul2/_086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_087_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_375_  (.A_N(net19),
    .B(\uut.mod_inv.sh1_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_088_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_376_  (.A0(\uut.mod_inv.mul_in1[0] ),
    .A1(net19),
    .S(\uut.mod_inv.sh1_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_089_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_377_  (.A(\uut.mod_inv.sh3_reg_1_1[0] ),
    .B_N(\uut.mod_inv.mul_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_090_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_378_  (.A0(\uut.mod_inv.mod_mul2/_088_ ),
    .A1(\uut.mod_inv.mod_mul2/_089_ ),
    .S(\uut.mod_inv.mod_mul2/_090_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_091_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_379_  (.A_N(net19),
    .B(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_092_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_380_  (.A0(\uut.mod_inv.mod_mul2/_189_ ),
    .A1(net19),
    .S(\uut.mod_inv.sh1_reg_1_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_093_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_381_  (.A(\uut.mod_inv.sh3_reg_1_1[2] ),
    .B_N(\uut.mod_inv.mul_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_094_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_382_  (.A0(\uut.mod_inv.mod_mul2/_092_ ),
    .A1(\uut.mod_inv.mod_mul2/_093_ ),
    .S(\uut.mod_inv.mod_mul2/_094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_095_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_383_  (.A(\uut.mod_inv.mod_mul2/_091_ ),
    .B(\uut.mod_inv.mod_mul2/_095_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_096_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_384_  (.A(\uut.mod_inv.mod_mul2/_087_ ),
    .B(\uut.mod_inv.mod_mul2/_096_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_097_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_385_  (.A_N(net15),
    .B(\uut.mod_inv.mod_mul2/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_098_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul2/_386_  (.A1(\uut.mod_inv.mod_mul2/_187_ ),
    .A2(\uut.mod_inv.mod_mul2/_020_ ),
    .B1_N(\uut.mod_inv.mod_mul2/_098_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_099_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_387_  (.A(\uut.mod_inv.sh3_reg_1_1[3] ),
    .B_N(\uut.mod_inv.mod_mul2/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_100_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_388_  (.A0(\uut.mod_inv.mod_mul2/_098_ ),
    .A1(\uut.mod_inv.mod_mul2/_099_ ),
    .S(\uut.mod_inv.mod_mul2/_100_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_101_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul2/_389_  (.A_N(\uut.mod_inv.sh3_reg_1_1[2] ),
    .B(\uut.mod_inv.mod_mul2/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_102_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_390_  (.A0(\uut.mod_inv.mod_mul2/_209_ ),
    .A1(\uut.mod_inv.sh3_reg_1_1[2] ),
    .S(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_103_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul2/_391_  (.A(net14),
    .B_N(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_104_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_392_  (.A0(\uut.mod_inv.mod_mul2/_102_ ),
    .A1(\uut.mod_inv.mod_mul2/_103_ ),
    .S(\uut.mod_inv.mod_mul2/_104_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_105_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_393_  (.A(\uut.mod_inv.mod_mul2/_002_ ),
    .B(\uut.mod_inv.mod_mul2/_105_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_106_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_394_  (.A(\uut.mod_inv.mod_mul2/_101_ ),
    .B(\uut.mod_inv.mod_mul2/_106_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_107_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_395_  (.A(\uut.mod_inv.mod_mul2/_197_ ),
    .B(\uut.mod_inv.mod_mul2/_213_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_108_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_396_  (.A(\uut.mod_inv.mod_mul2/_107_ ),
    .B(\uut.mod_inv.mod_mul2/_108_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_109_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_397_  (.A(\uut.mod_inv.mod_mul2/_097_ ),
    .B(\uut.mod_inv.mod_mul2/_109_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out2[2] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_398_  (.A(\uut.mod_inv.sh2_reg_1_1[2] ),
    .B(\uut.mod_inv.mod_mul2/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_110_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_399_  (.A(\uut.mod_inv.mod_mul2/_055_ ),
    .B(\uut.mod_inv.mod_mul2/_110_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_111_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_400_  (.A(net22),
    .B(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_112_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_401_  (.A1(net23),
    .A2(\uut.mod_inv.mod_mul2/_187_ ),
    .B1(\uut.mod_inv.mod_mul2/_020_ ),
    .B2(\uut.mod_inv.sh2_reg_1_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_113_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_402_  (.A(\uut.mod_inv.sh2_reg_1_1[3] ),
    .B(net23),
    .C(\uut.mod_inv.mod_mul2/_187_ ),
    .D(\uut.mod_inv.mod_mul2/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_114_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_403_  (.A(\uut.mod_inv.mod_mul2/_113_ ),
    .B(\uut.mod_inv.mod_mul2/_114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_115_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_404_  (.A(\uut.mod_inv.mod_mul2/_112_ ),
    .B(\uut.mod_inv.mod_mul2/_115_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_116_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_405_  (.A(\uut.mod_inv.mod_mul2/_111_ ),
    .B(\uut.mod_inv.mod_mul2/_116_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_117_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_406_  (.A(\uut.mod_inv.mod_mul2/_044_ ),
    .B(\uut.mod_inv.mod_mul2/_117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_118_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_407_  (.A(\uut.mod_inv.sh2_reg_1_1[2] ),
    .B(\uut.mod_inv.mod_mul2/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_119_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_408_  (.A(net26),
    .B(\uut.mod_inv.mod_mul2/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_120_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_409_  (.A(\uut.mod_inv.mod_mul2/_119_ ),
    .B(\uut.mod_inv.mod_mul2/_120_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_121_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_410_  (.A(\uut.mod_inv.mod_mul2/_036_ ),
    .B(\uut.mod_inv.mod_mul2/_121_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_122_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_411_  (.A(\uut.mod_inv.mod_mul2/_062_ ),
    .B(\uut.mod_inv.mod_mul2/_122_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_123_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul2/_412_  (.A1(net26),
    .A2(\uut.mod_inv.mod_mul2/_003_ ),
    .B1(\uut.mod_inv.mod_mul2/_189_ ),
    .B2(\uut.mod_inv.sh2_reg_1_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_124_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul2/_413_  (.A(\uut.mod_inv.sh2_reg_1_1[0] ),
    .B(net26),
    .C(\uut.mod_inv.mod_mul2/_003_ ),
    .D(\uut.mod_inv.mod_mul2/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_125_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_414_  (.A(\uut.mod_inv.mod_mul2/_124_ ),
    .B(\uut.mod_inv.mod_mul2/_125_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_126_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_415_  (.A(\uut.mod_inv.sh2_reg_1_1[0] ),
    .B(\uut.mod_inv.mod_mul2/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_127_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_416_  (.A(net23),
    .B(\uut.mod_inv.mod_mul2/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_128_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_417_  (.A(\uut.mod_inv.mod_mul2/_127_ ),
    .B(\uut.mod_inv.mod_mul2/_128_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_129_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_418_  (.A(\uut.mod_inv.mod_mul2/_126_ ),
    .B(\uut.mod_inv.mod_mul2/_129_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_130_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_419_  (.A(\uut.mod_inv.mod_mul2/_123_ ),
    .B(\uut.mod_inv.mod_mul2/_130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_131_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_420_  (.A(\uut.mod_inv.mod_mul2/_118_ ),
    .B(\uut.mod_inv.mod_mul2/_131_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out3[2] ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_421_  (.A(\uut.mod_inv.mod_mul2/_075_ ),
    .B(\uut.mod_inv.mod_mul2/_079_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_132_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul2/_422_  (.A(\uut.mod_inv.mod_mul2/_163_ ),
    .B(\uut.mod_inv.mod_mul2/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_133_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.mod_mul2/_423_  (.A(\uut.mod_inv.mod_mul2/_166_ ),
    .B(\uut.mod_inv.mod_mul2/_169_ ),
    .C(\uut.mod_inv.mod_mul2/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_134_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.mod_mul2/_424_  (.A(\uut.mod_inv.mod_mul2/_166_ ),
    .B(\uut.mod_inv.mod_mul2/_167_ ),
    .C(\uut.mod_inv.mod_mul2/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_135_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_425_  (.A(\uut.mod_inv.mod_mul2/_163_ ),
    .B(\uut.mod_inv.mod_mul2/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_136_ ));
 sky130_fd_sc_hd__a32o_1 \uut.mod_inv.mod_mul2/_426_  (.A1(\uut.mod_inv.mod_mul2/_133_ ),
    .A2(\uut.mod_inv.mod_mul2/_134_ ),
    .A3(\uut.mod_inv.mod_mul2/_135_ ),
    .B1(\uut.mod_inv.mod_mul2/_136_ ),
    .B2(\uut.mod_inv.mod_mul2/_170_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_137_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_427_  (.A(\uut.mod_inv.mod_mul2/_179_ ),
    .B(\uut.mod_inv.mod_mul2/_137_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_138_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.mod_mul2/_428_  (.A(\uut.mod_inv.mod_mul2/_162_ ),
    .B(\uut.mod_inv.mod_mul2/_166_ ),
    .C_N(\uut.mod_inv.mod_mul2/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_139_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul2/_429_  (.A(\uut.mod_inv.mod_mul2/_161_ ),
    .B(\uut.mod_inv.mod_mul2/_139_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_140_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.mod_mul2/_430_  (.A(\uut.mod_inv.mod_mul2/_160_ ),
    .B(\uut.mod_inv.mod_mul2/_166_ ),
    .C_N(\uut.mod_inv.mod_mul2/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_141_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_431_  (.A0(\uut.mod_inv.mod_mul2/_163_ ),
    .A1(\uut.mod_inv.mod_mul2/_070_ ),
    .S(\uut.mod_inv.mod_mul2/_141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_142_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul2/_432_  (.A0(\uut.mod_inv.mod_mul2/_140_ ),
    .A1(\uut.mod_inv.mod_mul2/_161_ ),
    .S(\uut.mod_inv.mod_mul2/_142_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_143_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_433_  (.A(\uut.mod_inv.mod_mul2/_138_ ),
    .B(\uut.mod_inv.mod_mul2/_143_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_144_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_434_  (.A(\uut.mod_inv.mod_mul2/_132_ ),
    .B(\uut.mod_inv.mod_mul2/_144_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out1[1] ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_435_  (.A(\uut.mod_inv.mod_mul2/_203_ ),
    .B(\uut.mod_inv.mod_mul2/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_145_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_436_  (.A(\uut.mod_inv.mod_mul2/_218_ ),
    .B(\uut.mod_inv.mod_mul2/_091_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_146_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_437_  (.A(\uut.mod_inv.mod_mul2/_107_ ),
    .B(\uut.mod_inv.mod_mul2/_146_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_147_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul2/_438_  (.A(\uut.mod_inv.mod_mul2/_145_ ),
    .B(\uut.mod_inv.mod_mul2/_147_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out2[1] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_439_  (.A(\uut.mod_inv.mod_mul2/_052_ ),
    .B(\uut.mod_inv.mod_mul2/_126_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_148_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_440_  (.A(\uut.mod_inv.mod_mul2/_041_ ),
    .B(\uut.mod_inv.mod_mul2/_117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_149_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul2/_441_  (.A(\uut.mod_inv.mod_mul2/_148_ ),
    .B(\uut.mod_inv.mod_mul2/_149_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out3[1] ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.mod_mul2/_442_  (.A1(\uut.mod_inv.mod_mul2/_162_ ),
    .A2(\uut.mod_inv.mod_mul2/_079_ ),
    .B1(\uut.mod_inv.mod_mul2/_076_ ),
    .B2(\uut.mod_inv.mod_mul2/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_150_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul2/_443_  (.A(\uut.mod_inv.mod_mul2/_159_ ),
    .B(\uut.mod_inv.mod_mul2/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_151_ ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.mod_mul2/_444_  (.A1(\uut.mod_inv.mod_mul2/_163_ ),
    .A2(\uut.mod_inv.mod_mul2/_151_ ),
    .B1(\uut.mod_inv.mod_mul2/_074_ ),
    .B2(\uut.mod_inv.mod_mul2/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_152_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_445_  (.A(\uut.mod_inv.mod_mul2/_150_ ),
    .B(\uut.mod_inv.mod_mul2/_152_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_153_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_446_  (.A(\uut.mod_inv.mod_mul2/_175_ ),
    .B(\uut.mod_inv.mod_mul2/_153_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_154_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_447_  (.A(\uut.mod_inv.mod_mul2/_172_ ),
    .B(\uut.mod_inv.mod_mul2/_154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out1[0] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul2/_448_  (.A(\uut.mod_inv.mod_mul2/_207_ ),
    .B(\uut.mod_inv.mod_mul2/_097_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul2/_155_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_449_  (.A(\uut.mod_inv.mod_mul2/_010_ ),
    .B(\uut.mod_inv.mod_mul2/_155_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out2[0] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_450_  (.A(\uut.mod_inv.mod_mul2/_058_ ),
    .B(\uut.mod_inv.mod_mul2/_130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_156_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_451_  (.A(\uut.mod_inv.mod_mul2/_066_ ),
    .B(\uut.mod_inv.mod_mul2/_122_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_157_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_452_  (.A(\uut.mod_inv.mod_mul2/_156_ ),
    .B(\uut.mod_inv.mod_mul2/_157_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2/_158_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul2/_453_  (.A(\uut.mod_inv.mod_mul2/_048_ ),
    .B(\uut.mod_inv.mod_mul2/_158_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul2_out3[0] ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul3/_221_  (.A(net17),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_159_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul3/_222_  (.A(\uut.mod_inv.sh3_reg_1_2[3] ),
    .B(\uut.mod_inv.sh2_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_160_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul3/_223_  (.A(\uut.mod_inv.mod_mul3/_159_ ),
    .B(\uut.mod_inv.mod_mul3/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_161_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul3/_224_  (.A(\uut.mod_inv.sh3_reg_1_2[2] ),
    .B(\uut.mod_inv.sh2_reg_1_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_162_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul3/_225_  (.A(net15),
    .B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_163_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_226_  (.A(\uut.mod_inv.mod_mul3/_162_ ),
    .B(\uut.mod_inv.mod_mul3/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_164_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_227_  (.A(\uut.mod_inv.mod_mul3/_161_ ),
    .B(\uut.mod_inv.mod_mul3/_164_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_165_ ));
 sky130_fd_sc_hd__xnor2_4 \uut.mod_inv.mod_mul3/_228_  (.A(\uut.mod_inv.mul_in3[3] ),
    .B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_166_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul3/_229_  (.A(\uut.mod_inv.sh3_reg_1_2[1] ),
    .B(\uut.mod_inv.sh2_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_167_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_230_  (.A(\uut.mod_inv.mod_mul3/_166_ ),
    .B(\uut.mod_inv.mod_mul3/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_168_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_231_  (.A(\uut.mod_inv.sh3_reg_1_2[1] ),
    .B(\uut.mod_inv.sh2_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_169_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_232_  (.A(\uut.mod_inv.mod_mul3/_166_ ),
    .B(\uut.mod_inv.mod_mul3/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_170_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_233_  (.A0(\uut.mod_inv.mod_mul3/_168_ ),
    .A1(\uut.mod_inv.mod_mul3/_170_ ),
    .S(\uut.mod_inv.mod_mul3/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_171_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_234_  (.A(\uut.mod_inv.mod_mul3/_165_ ),
    .B(\uut.mod_inv.mod_mul3/_171_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_172_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_235_  (.A(net19),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_173_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_236_  (.A(\uut.mod_inv.mod_mul3/_167_ ),
    .B(\uut.mod_inv.mod_mul3/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_174_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul3/_237_  (.A(\uut.mod_inv.mod_mul3/_169_ ),
    .B(\uut.mod_inv.mod_mul3/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_175_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_238_  (.A0(\uut.mod_inv.mod_mul3/_174_ ),
    .A1(\uut.mod_inv.mod_mul3/_175_ ),
    .S(\uut.mod_inv.mod_mul3/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_176_ ));
 sky130_fd_sc_hd__o22a_1 \uut.mod_inv.mod_mul3/_239_  (.A1(\uut.mod_inv.mod_mul3/_159_ ),
    .A2(\uut.mod_inv.mod_mul3/_162_ ),
    .B1(\uut.mod_inv.mod_mul3/_173_ ),
    .B2(\uut.mod_inv.mod_mul3/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_177_ ));
 sky130_fd_sc_hd__or4_1 \uut.mod_inv.mod_mul3/_240_  (.A(\uut.mod_inv.mod_mul3/_159_ ),
    .B(\uut.mod_inv.mod_mul3/_160_ ),
    .C(\uut.mod_inv.mod_mul3/_162_ ),
    .D(\uut.mod_inv.mod_mul3/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_178_ ));
 sky130_fd_sc_hd__nor2b_1 \uut.mod_inv.mod_mul3/_241_  (.A(\uut.mod_inv.mod_mul3/_177_ ),
    .B_N(\uut.mod_inv.mod_mul3/_178_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_179_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_242_  (.A(\uut.mod_inv.mod_mul3/_159_ ),
    .B(\uut.mod_inv.mod_mul3/_167_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_180_ ));
 sky130_fd_sc_hd__xor2_2 \uut.mod_inv.mod_mul3/_243_  (.A(\uut.mod_inv.sh3_reg_1_2[0] ),
    .B(\uut.mod_inv.sh2_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_181_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_244_  (.A0(\uut.mod_inv.mod_mul3/_167_ ),
    .A1(\uut.mod_inv.mod_mul3/_181_ ),
    .S(\uut.mod_inv.mod_mul3/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_182_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_245_  (.A(\uut.mod_inv.mod_mul3/_166_ ),
    .B(\uut.mod_inv.mod_mul3/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_183_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_246_  (.A0(\uut.mod_inv.mod_mul3/_180_ ),
    .A1(\uut.mod_inv.mod_mul3/_182_ ),
    .S(\uut.mod_inv.mod_mul3/_183_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_184_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_247_  (.A(\uut.mod_inv.mod_mul3/_179_ ),
    .B(\uut.mod_inv.mod_mul3/_184_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_185_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_248_  (.A(\uut.mod_inv.mod_mul3/_176_ ),
    .B(\uut.mod_inv.mod_mul3/_185_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_186_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_249_  (.A(\uut.mod_inv.mod_mul3/_172_ ),
    .B(\uut.mod_inv.mod_mul3/_186_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out1[3] ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_250_  (.A(\uut.mod_inv.sh1_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_187_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_251_  (.A_N(net19),
    .B(\uut.mod_inv.mod_mul3/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_188_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_252_  (.A(\uut.mod_inv.mul_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_189_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul3/_253_  (.A1(\uut.mod_inv.mod_mul3/_187_ ),
    .A2(\uut.mod_inv.mod_mul3/_189_ ),
    .B1_N(\uut.mod_inv.mod_mul3/_188_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_190_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_254_  (.A(\uut.mod_inv.sh3_reg_1_2[3] ),
    .B_N(\uut.mod_inv.mod_mul3/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_191_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_255_  (.A0(\uut.mod_inv.mod_mul3/_188_ ),
    .A1(\uut.mod_inv.mod_mul3/_190_ ),
    .S(\uut.mod_inv.mod_mul3/_191_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_192_ ));
 sky130_fd_sc_hd__clkbuf_4 \uut.mod_inv.mod_mul3/_256_  (.A(\uut.mod_inv.sh1_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_193_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_257_  (.A_N(net18),
    .B(\uut.mod_inv.mod_mul3/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_194_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_258_  (.A0(net20),
    .A1(net18),
    .S(\uut.mod_inv.sh1_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_195_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_259_  (.A(\uut.mod_inv.sh3_reg_1_2[1] ),
    .B_N(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_196_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul3/_260_  (.A0(\uut.mod_inv.mod_mul3/_194_ ),
    .A1(\uut.mod_inv.mod_mul3/_195_ ),
    .S(\uut.mod_inv.mod_mul3/_196_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_197_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_261_  (.A_N(net18),
    .B(\uut.mod_inv.sh1_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_198_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_262_  (.A0(net20),
    .A1(net18),
    .S(\uut.mod_inv.sh1_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_199_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_263_  (.A(\uut.mod_inv.sh3_reg_1_2[3] ),
    .B_N(\uut.mod_inv.mul_in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_200_ ));
 sky130_fd_sc_hd__mux2_2 \uut.mod_inv.mod_mul3/_264_  (.A0(\uut.mod_inv.mod_mul3/_198_ ),
    .A1(\uut.mod_inv.mod_mul3/_199_ ),
    .S(\uut.mod_inv.mod_mul3/_200_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_201_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_265_  (.A(\uut.mod_inv.mod_mul3/_197_ ),
    .B(\uut.mod_inv.mod_mul3/_201_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_202_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_266_  (.A(\uut.mod_inv.mod_mul3/_192_ ),
    .B(\uut.mod_inv.mod_mul3/_202_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_203_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_267_  (.A_N(net19),
    .B(\uut.mod_inv.mod_mul3/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_204_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul3/_268_  (.A1(\uut.mod_inv.mod_mul3/_193_ ),
    .A2(\uut.mod_inv.mod_mul3/_189_ ),
    .B1_N(\uut.mod_inv.mod_mul3/_204_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_205_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_269_  (.A(\uut.mod_inv.sh3_reg_1_2[1] ),
    .B_N(\uut.mod_inv.mod_mul3/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_206_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_270_  (.A0(\uut.mod_inv.mod_mul3/_204_ ),
    .A1(\uut.mod_inv.mod_mul3/_205_ ),
    .S(\uut.mod_inv.mod_mul3/_206_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_207_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_271_  (.A(\uut.mod_inv.mod_mul3/_203_ ),
    .B(\uut.mod_inv.mod_mul3/_207_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_208_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_272_  (.A(\uut.mod_inv.sh1_reg_1_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_209_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_273_  (.A_N(net16),
    .B(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_210_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_274_  (.A0(\uut.mod_inv.mul_in1[2] ),
    .A1(net16),
    .S(\uut.mod_inv.sh1_reg_1_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_211_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_275_  (.A(\uut.mod_inv.sh3_reg_1_2[2] ),
    .B_N(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_212_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_276_  (.A0(\uut.mod_inv.mod_mul3/_210_ ),
    .A1(\uut.mod_inv.mod_mul3/_211_ ),
    .S(\uut.mod_inv.mod_mul3/_212_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_213_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_277_  (.A_N(net14),
    .B(\uut.mod_inv.sh1_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_214_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_278_  (.A(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_215_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_279_  (.A0(\uut.mod_inv.mod_mul3/_215_ ),
    .A1(net14),
    .S(\uut.mod_inv.sh1_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_216_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_280_  (.A(\uut.mod_inv.sh3_reg_1_2[3] ),
    .B_N(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_217_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_281_  (.A0(\uut.mod_inv.mod_mul3/_214_ ),
    .A1(\uut.mod_inv.mod_mul3/_216_ ),
    .S(\uut.mod_inv.mod_mul3/_217_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_218_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_282_  (.A(\uut.mod_inv.mod_mul3/_213_ ),
    .B(\uut.mod_inv.mod_mul3/_218_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_219_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_283_  (.A_N(\uut.mod_inv.sh3_reg_1_2[1] ),
    .B(\uut.mod_inv.mod_mul3/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_220_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_284_  (.A0(\uut.mod_inv.sh1_reg_1_2[1] ),
    .A1(\uut.mod_inv.sh3_reg_1_2[1] ),
    .S(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_000_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_285_  (.A(net14),
    .B_N(\uut.mod_inv.sh1_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_001_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_286_  (.A0(\uut.mod_inv.mod_mul3/_220_ ),
    .A1(\uut.mod_inv.mod_mul3/_000_ ),
    .S(\uut.mod_inv.mod_mul3/_001_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_002_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_287_  (.A(\uut.mod_inv.sh1_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_003_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_288_  (.A_N(net18),
    .B(\uut.mod_inv.mod_mul3/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_004_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_289_  (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_005_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_290_  (.A0(\uut.mod_inv.mod_mul3/_005_ ),
    .A1(net18),
    .S(\uut.mod_inv.sh1_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_006_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_291_  (.A(\uut.mod_inv.sh3_reg_1_2[0] ),
    .B_N(\uut.mod_inv.mod_mul3/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_007_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_292_  (.A0(\uut.mod_inv.mod_mul3/_004_ ),
    .A1(\uut.mod_inv.mod_mul3/_006_ ),
    .S(\uut.mod_inv.mod_mul3/_007_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_008_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_293_  (.A(\uut.mod_inv.mod_mul3/_002_ ),
    .B(\uut.mod_inv.mod_mul3/_008_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_009_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_294_  (.A(\uut.mod_inv.mod_mul3/_219_ ),
    .B(\uut.mod_inv.mod_mul3/_009_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_010_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_295_  (.A_N(\uut.mod_inv.sh3_reg_1_2[0] ),
    .B(\uut.mod_inv.mod_mul3/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_011_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul3/_296_  (.A1(\uut.mod_inv.mod_mul3/_215_ ),
    .A2(\uut.mod_inv.mod_mul3/_003_ ),
    .B1_N(\uut.mod_inv.mod_mul3/_011_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_012_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_297_  (.A(net14),
    .B_N(\uut.mod_inv.mod_mul3/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_013_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_298_  (.A0(\uut.mod_inv.mod_mul3/_011_ ),
    .A1(\uut.mod_inv.mod_mul3/_012_ ),
    .S(\uut.mod_inv.mod_mul3/_013_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_014_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_299_  (.A_N(net18),
    .B(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_015_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_300_  (.A0(\uut.mod_inv.mod_mul3/_005_ ),
    .A1(net18),
    .S(\uut.mod_inv.sh1_reg_1_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_016_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_301_  (.A(\uut.mod_inv.sh3_reg_1_2[2] ),
    .B_N(\uut.mod_inv.mul_in1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_017_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_302_  (.A0(\uut.mod_inv.mod_mul3/_015_ ),
    .A1(\uut.mod_inv.mod_mul3/_016_ ),
    .S(\uut.mod_inv.mod_mul3/_017_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_018_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_303_  (.A_N(net16),
    .B(\uut.mod_inv.mod_mul3/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_019_ ));
 sky130_fd_sc_hd__buf_2 \uut.mod_inv.mod_mul3/_304_  (.A(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_020_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_305_  (.A0(\uut.mod_inv.mod_mul3/_020_ ),
    .A1(net16),
    .S(\uut.mod_inv.sh1_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_021_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_306_  (.A(\uut.mod_inv.sh3_reg_1_2[1] ),
    .B_N(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_022_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_307_  (.A0(\uut.mod_inv.mod_mul3/_019_ ),
    .A1(\uut.mod_inv.mod_mul3/_021_ ),
    .S(\uut.mod_inv.mod_mul3/_022_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_023_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_308_  (.A(\uut.mod_inv.mod_mul3/_018_ ),
    .B(\uut.mod_inv.mod_mul3/_023_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_024_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_309_  (.A(\uut.mod_inv.mod_mul3/_014_ ),
    .B(\uut.mod_inv.mod_mul3/_024_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_025_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_310_  (.A(\uut.mod_inv.mod_mul3/_010_ ),
    .B(\uut.mod_inv.mod_mul3/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_026_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_311_  (.A(\uut.mod_inv.mod_mul3/_208_ ),
    .B(\uut.mod_inv.mod_mul3/_026_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out2[3] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_312_  (.A(net25),
    .B(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_027_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_313_  (.A(\uut.mod_inv.sh2_reg_1_2[2] ),
    .B(\uut.mod_inv.mod_mul3/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_028_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_314_  (.A(\uut.mod_inv.mod_mul3/_027_ ),
    .B(\uut.mod_inv.mod_mul3/_028_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_029_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_315_  (.A(net26),
    .B(\uut.mod_inv.mod_mul3/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_030_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_316_  (.A(\uut.mod_inv.sh2_reg_1_2[3] ),
    .B(\uut.mod_inv.mod_mul3/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_031_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_317_  (.A(\uut.mod_inv.mod_mul3/_030_ ),
    .B(\uut.mod_inv.mod_mul3/_031_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_032_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_318_  (.A(\uut.mod_inv.mod_mul3/_029_ ),
    .B(\uut.mod_inv.mod_mul3/_032_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_033_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_319_  (.A1(net25),
    .A2(\uut.mod_inv.mod_mul3/_187_ ),
    .B1(\uut.mod_inv.mod_mul3/_005_ ),
    .B2(\uut.mod_inv.sh2_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_034_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_320_  (.A(\uut.mod_inv.sh2_reg_1_2[3] ),
    .B(net25),
    .C(\uut.mod_inv.mod_mul3/_187_ ),
    .D(\uut.mod_inv.mod_mul3/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_035_ ));
 sky130_fd_sc_hd__nor2_2 \uut.mod_inv.mod_mul3/_321_  (.A(\uut.mod_inv.mod_mul3/_034_ ),
    .B(\uut.mod_inv.mod_mul3/_035_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_036_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_322_  (.A(\uut.mod_inv.inv_out3_xor[2] ),
    .B(\uut.mod_inv.mod_mul3/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_037_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_323_  (.A(\uut.mod_inv.sh2_reg_1_2[1] ),
    .B(\uut.mod_inv.mod_mul3/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_038_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_324_  (.A(\uut.mod_inv.mod_mul3/_037_ ),
    .B(\uut.mod_inv.mod_mul3/_038_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_039_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_325_  (.A(\uut.mod_inv.mod_mul3/_036_ ),
    .B(\uut.mod_inv.mod_mul3/_039_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_040_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_326_  (.A(\uut.mod_inv.mod_mul3/_033_ ),
    .B(\uut.mod_inv.mod_mul3/_040_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_041_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_327_  (.A1(\uut.mod_inv.sh2_reg_1_2[1] ),
    .A2(\uut.mod_inv.mod_mul3/_215_ ),
    .B1(\uut.mod_inv.mod_mul3/_193_ ),
    .B2(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_042_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_328_  (.A(net22),
    .B(\uut.mod_inv.sh2_reg_1_2[1] ),
    .C(\uut.mod_inv.mod_mul3/_215_ ),
    .D(\uut.mod_inv.mod_mul3/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_043_ ));
 sky130_fd_sc_hd__nor2_2 \uut.mod_inv.mod_mul3/_329_  (.A(\uut.mod_inv.mod_mul3/_042_ ),
    .B(\uut.mod_inv.mod_mul3/_043_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_044_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_330_  (.A(\uut.mod_inv.sh2_reg_1_2[3] ),
    .B(\uut.mod_inv.mod_mul3/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_045_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_331_  (.A(\uut.mod_inv.inv_out3_xor[3] ),
    .B(\uut.mod_inv.mod_mul3/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_046_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_332_  (.A(\uut.mod_inv.mod_mul3/_045_ ),
    .B(\uut.mod_inv.mod_mul3/_046_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_047_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_333_  (.A(\uut.mod_inv.mod_mul3/_044_ ),
    .B(\uut.mod_inv.mod_mul3/_047_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_048_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_334_  (.A(\uut.mod_inv.sh2_reg_1_2[0] ),
    .B(\uut.mod_inv.mod_mul3/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_049_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_335_  (.A(\uut.mod_inv.inv_out3_xor[3] ),
    .B(\uut.mod_inv.mod_mul3/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_050_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_336_  (.A(\uut.mod_inv.mod_mul3/_049_ ),
    .B(\uut.mod_inv.mod_mul3/_050_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_051_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_337_  (.A(\uut.mod_inv.mod_mul3/_048_ ),
    .B(\uut.mod_inv.mod_mul3/_051_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_052_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_338_  (.A1(net24),
    .A2(\uut.mod_inv.mod_mul3/_193_ ),
    .B1(\uut.mod_inv.mod_mul3/_005_ ),
    .B2(\uut.mod_inv.sh2_reg_1_2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_053_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_339_  (.A(\uut.mod_inv.sh2_reg_1_2[1] ),
    .B(net25),
    .C(\uut.mod_inv.mod_mul3/_193_ ),
    .D(\uut.mod_inv.mod_mul3/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_054_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_340_  (.A(\uut.mod_inv.mod_mul3/_053_ ),
    .B(\uut.mod_inv.mod_mul3/_054_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_055_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_341_  (.A1(net25),
    .A2(\uut.mod_inv.mod_mul3/_003_ ),
    .B1(\uut.mod_inv.mod_mul3/_005_ ),
    .B2(\uut.mod_inv.sh2_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_056_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_342_  (.A(\uut.mod_inv.sh2_reg_1_2[0] ),
    .B(net25),
    .C(\uut.mod_inv.mod_mul3/_003_ ),
    .D(\uut.mod_inv.mod_mul3/_005_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_057_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_343_  (.A(\uut.mod_inv.mod_mul3/_056_ ),
    .B(\uut.mod_inv.mod_mul3/_057_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_058_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_344_  (.A(\uut.mod_inv.mod_mul3/_055_ ),
    .B(\uut.mod_inv.mod_mul3/_058_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_059_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_345_  (.A1(\uut.mod_inv.inv_out3_xor[2] ),
    .A2(\uut.mod_inv.mod_mul3/_209_ ),
    .B1(\uut.mod_inv.mod_mul3/_020_ ),
    .B2(\uut.mod_inv.sh2_reg_1_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_060_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_346_  (.A(\uut.mod_inv.sh2_reg_1_2[2] ),
    .B(net23),
    .C(\uut.mod_inv.mod_mul3/_209_ ),
    .D(\uut.mod_inv.mod_mul3/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_061_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_347_  (.A(\uut.mod_inv.mod_mul3/_060_ ),
    .B(\uut.mod_inv.mod_mul3/_061_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_062_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_348_  (.A(\uut.mod_inv.sh2_reg_1_2[1] ),
    .B(\uut.mod_inv.mod_mul3/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_063_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_349_  (.A(net26),
    .B(\uut.mod_inv.mod_mul3/_193_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_064_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_350_  (.A(\uut.mod_inv.mod_mul3/_063_ ),
    .B(\uut.mod_inv.mod_mul3/_064_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_065_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_351_  (.A(\uut.mod_inv.mod_mul3/_062_ ),
    .B(\uut.mod_inv.mod_mul3/_065_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_066_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_352_  (.A(\uut.mod_inv.mod_mul3/_059_ ),
    .B(\uut.mod_inv.mod_mul3/_066_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_067_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_353_  (.A(\uut.mod_inv.mod_mul3/_052_ ),
    .B(\uut.mod_inv.mod_mul3/_067_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_068_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_354_  (.A(\uut.mod_inv.mod_mul3/_041_ ),
    .B(\uut.mod_inv.mod_mul3/_068_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out3[3] ));
 sky130_fd_sc_hd__a21bo_1 \uut.mod_inv.mod_mul3/_355_  (.A1(\uut.mod_inv.mod_mul3/_160_ ),
    .A2(\uut.mod_inv.mod_mul3/_164_ ),
    .B1_N(\uut.mod_inv.mod_mul3/_161_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_069_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_356_  (.A(\uut.mod_inv.mod_mul3/_160_ ),
    .B(\uut.mod_inv.mod_mul3/_163_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_070_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_357_  (.A(\uut.mod_inv.mod_mul3/_162_ ),
    .B(\uut.mod_inv.mod_mul3/_070_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_071_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_358_  (.A0(\uut.mod_inv.mod_mul3/_159_ ),
    .A1(\uut.mod_inv.mod_mul3/_069_ ),
    .S(\uut.mod_inv.mod_mul3/_071_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_072_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_359_  (.A(\uut.mod_inv.sh3_reg_1_2[0] ),
    .B(\uut.mod_inv.sh2_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_073_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_360_  (.A(\uut.mod_inv.mod_mul3/_163_ ),
    .B(\uut.mod_inv.mod_mul3/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_074_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul3/_361_  (.A(\uut.mod_inv.mod_mul3/_159_ ),
    .B(\uut.mod_inv.mod_mul3/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_075_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_362_  (.A(\uut.mod_inv.mod_mul3/_162_ ),
    .B(\uut.mod_inv.mod_mul3/_173_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_076_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_363_  (.A(\uut.mod_inv.mod_mul3/_075_ ),
    .B(\uut.mod_inv.mod_mul3/_076_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_364_  (.A(\uut.mod_inv.mod_mul3/_074_ ),
    .B(\uut.mod_inv.mod_mul3/_077_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_078_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_365_  (.A(\uut.mod_inv.mod_mul3/_173_ ),
    .B(\uut.mod_inv.mod_mul3/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_079_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_366_  (.A0(\uut.mod_inv.mod_mul3/_168_ ),
    .A1(\uut.mod_inv.mod_mul3/_170_ ),
    .S(\uut.mod_inv.mod_mul3/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_080_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_367_  (.A(\uut.mod_inv.mod_mul3/_079_ ),
    .B(\uut.mod_inv.mod_mul3/_080_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_081_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_368_  (.A(\uut.mod_inv.mod_mul3/_078_ ),
    .B(\uut.mod_inv.mod_mul3/_081_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_082_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_369_  (.A(\uut.mod_inv.mod_mul3/_072_ ),
    .B(\uut.mod_inv.mod_mul3/_082_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out1[2] ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_370_  (.A_N(net16),
    .B(\uut.mod_inv.mod_mul3/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_083_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_371_  (.A0(\uut.mod_inv.mod_mul3/_020_ ),
    .A1(net15),
    .S(\uut.mod_inv.sh1_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_084_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_372_  (.A(\uut.mod_inv.sh3_reg_1_2[0] ),
    .B_N(\uut.mod_inv.mul_in1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_085_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_373_  (.A0(\uut.mod_inv.mod_mul3/_083_ ),
    .A1(\uut.mod_inv.mod_mul3/_084_ ),
    .S(\uut.mod_inv.mod_mul3/_085_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_086_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_374_  (.A(\uut.mod_inv.mod_mul3/_201_ ),
    .B(\uut.mod_inv.mod_mul3/_086_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_087_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_375_  (.A_N(\uut.mod_inv.mul_in3[0] ),
    .B(\uut.mod_inv.sh1_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_088_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_376_  (.A0(\uut.mod_inv.mul_in1[0] ),
    .A1(\uut.mod_inv.mul_in3[0] ),
    .S(\uut.mod_inv.sh1_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_089_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_377_  (.A(\uut.mod_inv.sh3_reg_1_2[0] ),
    .B_N(\uut.mod_inv.mul_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_090_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_378_  (.A0(\uut.mod_inv.mod_mul3/_088_ ),
    .A1(\uut.mod_inv.mod_mul3/_089_ ),
    .S(\uut.mod_inv.mod_mul3/_090_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_091_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_379_  (.A_N(\uut.mod_inv.mul_in3[0] ),
    .B(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_092_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_380_  (.A0(\uut.mod_inv.mod_mul3/_189_ ),
    .A1(\uut.mod_inv.mul_in3[0] ),
    .S(\uut.mod_inv.sh1_reg_1_2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_093_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_381_  (.A(\uut.mod_inv.sh3_reg_1_2[2] ),
    .B_N(\uut.mod_inv.mul_in1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_094_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_382_  (.A0(\uut.mod_inv.mod_mul3/_092_ ),
    .A1(\uut.mod_inv.mod_mul3/_093_ ),
    .S(\uut.mod_inv.mod_mul3/_094_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_095_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_383_  (.A(\uut.mod_inv.mod_mul3/_091_ ),
    .B(\uut.mod_inv.mod_mul3/_095_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_096_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_384_  (.A(\uut.mod_inv.mod_mul3/_087_ ),
    .B(\uut.mod_inv.mod_mul3/_096_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_097_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_385_  (.A_N(net16),
    .B(\uut.mod_inv.mod_mul3/_187_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_098_ ));
 sky130_fd_sc_hd__o21ba_1 \uut.mod_inv.mod_mul3/_386_  (.A1(\uut.mod_inv.mod_mul3/_187_ ),
    .A2(\uut.mod_inv.mod_mul3/_020_ ),
    .B1_N(\uut.mod_inv.mod_mul3/_098_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_099_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_387_  (.A(\uut.mod_inv.sh3_reg_1_2[3] ),
    .B_N(\uut.mod_inv.mod_mul3/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_100_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_388_  (.A0(\uut.mod_inv.mod_mul3/_098_ ),
    .A1(\uut.mod_inv.mod_mul3/_099_ ),
    .S(\uut.mod_inv.mod_mul3/_100_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_101_ ));
 sky130_fd_sc_hd__and2b_1 \uut.mod_inv.mod_mul3/_389_  (.A_N(\uut.mod_inv.sh3_reg_1_2[2] ),
    .B(\uut.mod_inv.mod_mul3/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_102_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_390_  (.A0(\uut.mod_inv.mod_mul3/_209_ ),
    .A1(\uut.mod_inv.sh3_reg_1_2[2] ),
    .S(\uut.mod_inv.mul_in1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_103_ ));
 sky130_fd_sc_hd__or2b_1 \uut.mod_inv.mod_mul3/_391_  (.A(\uut.mod_inv.mul_in3[3] ),
    .B_N(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_104_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_392_  (.A0(\uut.mod_inv.mod_mul3/_102_ ),
    .A1(\uut.mod_inv.mod_mul3/_103_ ),
    .S(\uut.mod_inv.mod_mul3/_104_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_105_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_393_  (.A(\uut.mod_inv.mod_mul3/_002_ ),
    .B(\uut.mod_inv.mod_mul3/_105_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_106_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_394_  (.A(\uut.mod_inv.mod_mul3/_101_ ),
    .B(\uut.mod_inv.mod_mul3/_106_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_107_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_395_  (.A(\uut.mod_inv.mod_mul3/_197_ ),
    .B(\uut.mod_inv.mod_mul3/_213_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_108_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_396_  (.A(\uut.mod_inv.mod_mul3/_107_ ),
    .B(\uut.mod_inv.mod_mul3/_108_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_109_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_397_  (.A(\uut.mod_inv.mod_mul3/_097_ ),
    .B(\uut.mod_inv.mod_mul3/_109_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out2[2] ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_398_  (.A(\uut.mod_inv.sh2_reg_1_2[2] ),
    .B(\uut.mod_inv.mod_mul3/_215_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_110_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_399_  (.A(\uut.mod_inv.mod_mul3/_055_ ),
    .B(\uut.mod_inv.mod_mul3/_110_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_111_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_400_  (.A(net22),
    .B(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_112_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_401_  (.A1(\uut.mod_inv.inv_out3_xor[2] ),
    .A2(\uut.mod_inv.mod_mul3/_187_ ),
    .B1(\uut.mod_inv.mod_mul3/_020_ ),
    .B2(\uut.mod_inv.sh2_reg_1_2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_113_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_402_  (.A(\uut.mod_inv.sh2_reg_1_2[3] ),
    .B(\uut.mod_inv.inv_out3_xor[2] ),
    .C(\uut.mod_inv.mod_mul3/_187_ ),
    .D(\uut.mod_inv.mod_mul3/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_114_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_403_  (.A(\uut.mod_inv.mod_mul3/_113_ ),
    .B(\uut.mod_inv.mod_mul3/_114_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_115_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_404_  (.A(\uut.mod_inv.mod_mul3/_112_ ),
    .B(\uut.mod_inv.mod_mul3/_115_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_116_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_405_  (.A(\uut.mod_inv.mod_mul3/_111_ ),
    .B(\uut.mod_inv.mod_mul3/_116_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_117_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_406_  (.A(\uut.mod_inv.mod_mul3/_044_ ),
    .B(\uut.mod_inv.mod_mul3/_117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_118_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_407_  (.A(\uut.mod_inv.sh2_reg_1_2[2] ),
    .B(\uut.mod_inv.mod_mul3/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_119_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_408_  (.A(net26),
    .B(\uut.mod_inv.mod_mul3/_209_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_120_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_409_  (.A(\uut.mod_inv.mod_mul3/_119_ ),
    .B(\uut.mod_inv.mod_mul3/_120_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_121_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_410_  (.A(\uut.mod_inv.mod_mul3/_036_ ),
    .B(\uut.mod_inv.mod_mul3/_121_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_122_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_411_  (.A(\uut.mod_inv.mod_mul3/_062_ ),
    .B(\uut.mod_inv.mod_mul3/_122_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_123_ ));
 sky130_fd_sc_hd__a22oi_1 \uut.mod_inv.mod_mul3/_412_  (.A1(\uut.mod_inv.inv_out3_xor[0] ),
    .A2(\uut.mod_inv.mod_mul3/_003_ ),
    .B1(\uut.mod_inv.mod_mul3/_189_ ),
    .B2(\uut.mod_inv.sh2_reg_1_2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_124_ ));
 sky130_fd_sc_hd__and4_1 \uut.mod_inv.mod_mul3/_413_  (.A(\uut.mod_inv.sh2_reg_1_2[0] ),
    .B(\uut.mod_inv.inv_out3_xor[0] ),
    .C(\uut.mod_inv.mod_mul3/_003_ ),
    .D(\uut.mod_inv.mod_mul3/_189_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_125_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_414_  (.A(\uut.mod_inv.mod_mul3/_124_ ),
    .B(\uut.mod_inv.mod_mul3/_125_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_126_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_415_  (.A(\uut.mod_inv.sh2_reg_1_2[0] ),
    .B(\uut.mod_inv.mod_mul3/_020_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_127_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_416_  (.A(net23),
    .B(\uut.mod_inv.mod_mul3/_003_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_128_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_417_  (.A(\uut.mod_inv.mod_mul3/_127_ ),
    .B(\uut.mod_inv.mod_mul3/_128_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_129_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_418_  (.A(\uut.mod_inv.mod_mul3/_126_ ),
    .B(\uut.mod_inv.mod_mul3/_129_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_130_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_419_  (.A(\uut.mod_inv.mod_mul3/_123_ ),
    .B(\uut.mod_inv.mod_mul3/_130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_131_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_420_  (.A(\uut.mod_inv.mod_mul3/_118_ ),
    .B(\uut.mod_inv.mod_mul3/_131_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out3[2] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_421_  (.A(\uut.mod_inv.mod_mul3/_075_ ),
    .B(\uut.mod_inv.mod_mul3/_079_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_132_ ));
 sky130_fd_sc_hd__or2_1 \uut.mod_inv.mod_mul3/_422_  (.A(\uut.mod_inv.mod_mul3/_163_ ),
    .B(\uut.mod_inv.mod_mul3/_169_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_133_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.mod_mul3/_423_  (.A(\uut.mod_inv.mod_mul3/_166_ ),
    .B(\uut.mod_inv.mod_mul3/_169_ ),
    .C(\uut.mod_inv.mod_mul3/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_134_ ));
 sky130_fd_sc_hd__or3_1 \uut.mod_inv.mod_mul3/_424_  (.A(\uut.mod_inv.mod_mul3/_166_ ),
    .B(\uut.mod_inv.mod_mul3/_167_ ),
    .C(\uut.mod_inv.mod_mul3/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_135_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_425_  (.A(\uut.mod_inv.mod_mul3/_163_ ),
    .B(\uut.mod_inv.mod_mul3/_181_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_136_ ));
 sky130_fd_sc_hd__a32o_1 \uut.mod_inv.mod_mul3/_426_  (.A1(\uut.mod_inv.mod_mul3/_133_ ),
    .A2(\uut.mod_inv.mod_mul3/_134_ ),
    .A3(\uut.mod_inv.mod_mul3/_135_ ),
    .B1(\uut.mod_inv.mod_mul3/_136_ ),
    .B2(\uut.mod_inv.mod_mul3/_170_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_137_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_427_  (.A(\uut.mod_inv.mod_mul3/_179_ ),
    .B(\uut.mod_inv.mod_mul3/_137_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_138_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.mod_mul3/_428_  (.A(\uut.mod_inv.mod_mul3/_162_ ),
    .B(\uut.mod_inv.mod_mul3/_166_ ),
    .C_N(\uut.mod_inv.mod_mul3/_160_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_139_ ));
 sky130_fd_sc_hd__nand2_1 \uut.mod_inv.mod_mul3/_429_  (.A(\uut.mod_inv.mod_mul3/_161_ ),
    .B(\uut.mod_inv.mod_mul3/_139_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_140_ ));
 sky130_fd_sc_hd__or3b_1 \uut.mod_inv.mod_mul3/_430_  (.A(\uut.mod_inv.mod_mul3/_160_ ),
    .B(\uut.mod_inv.mod_mul3/_166_ ),
    .C_N(\uut.mod_inv.mod_mul3/_162_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_141_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_431_  (.A0(\uut.mod_inv.mod_mul3/_163_ ),
    .A1(\uut.mod_inv.mod_mul3/_070_ ),
    .S(\uut.mod_inv.mod_mul3/_141_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_142_ ));
 sky130_fd_sc_hd__mux2_1 \uut.mod_inv.mod_mul3/_432_  (.A0(\uut.mod_inv.mod_mul3/_140_ ),
    .A1(\uut.mod_inv.mod_mul3/_161_ ),
    .S(\uut.mod_inv.mod_mul3/_142_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_143_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_433_  (.A(\uut.mod_inv.mod_mul3/_138_ ),
    .B(\uut.mod_inv.mod_mul3/_143_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_144_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_434_  (.A(\uut.mod_inv.mod_mul3/_132_ ),
    .B(\uut.mod_inv.mod_mul3/_144_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out1[1] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_435_  (.A(\uut.mod_inv.mod_mul3/_203_ ),
    .B(\uut.mod_inv.mod_mul3/_025_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_145_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_436_  (.A(\uut.mod_inv.mod_mul3/_218_ ),
    .B(\uut.mod_inv.mod_mul3/_091_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_146_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_437_  (.A(\uut.mod_inv.mod_mul3/_107_ ),
    .B(\uut.mod_inv.mod_mul3/_146_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_147_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_438_  (.A(\uut.mod_inv.mod_mul3/_145_ ),
    .B(\uut.mod_inv.mod_mul3/_147_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out2[1] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_439_  (.A(\uut.mod_inv.mod_mul3/_052_ ),
    .B(\uut.mod_inv.mod_mul3/_126_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_148_ ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_440_  (.A(\uut.mod_inv.mod_mul3/_041_ ),
    .B(\uut.mod_inv.mod_mul3/_117_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_149_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_441_  (.A(\uut.mod_inv.mod_mul3/_148_ ),
    .B(\uut.mod_inv.mod_mul3/_149_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out3[1] ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.mod_mul3/_442_  (.A1(\uut.mod_inv.mod_mul3/_162_ ),
    .A2(\uut.mod_inv.mod_mul3/_079_ ),
    .B1(\uut.mod_inv.mod_mul3/_076_ ),
    .B2(\uut.mod_inv.mod_mul3/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_150_ ));
 sky130_fd_sc_hd__nor2_1 \uut.mod_inv.mod_mul3/_443_  (.A(\uut.mod_inv.mod_mul3/_159_ ),
    .B(\uut.mod_inv.mod_mul3/_073_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_151_ ));
 sky130_fd_sc_hd__a22o_1 \uut.mod_inv.mod_mul3/_444_  (.A1(\uut.mod_inv.mod_mul3/_163_ ),
    .A2(\uut.mod_inv.mod_mul3/_151_ ),
    .B1(\uut.mod_inv.mod_mul3/_074_ ),
    .B2(\uut.mod_inv.mod_mul3/_159_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_152_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_445_  (.A(\uut.mod_inv.mod_mul3/_150_ ),
    .B(\uut.mod_inv.mod_mul3/_152_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_153_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_446_  (.A(\uut.mod_inv.mod_mul3/_175_ ),
    .B(\uut.mod_inv.mod_mul3/_153_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_154_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_447_  (.A(\uut.mod_inv.mod_mul3/_172_ ),
    .B(\uut.mod_inv.mod_mul3/_154_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out1[0] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.mod_mul3/_448_  (.A(\uut.mod_inv.mod_mul3/_207_ ),
    .B(\uut.mod_inv.mod_mul3/_097_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.mod_mul3/_155_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_449_  (.A(\uut.mod_inv.mod_mul3/_010_ ),
    .B(\uut.mod_inv.mod_mul3/_155_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out2[0] ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_450_  (.A(\uut.mod_inv.mod_mul3/_058_ ),
    .B(\uut.mod_inv.mod_mul3/_130_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_156_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_451_  (.A(\uut.mod_inv.mod_mul3/_066_ ),
    .B(\uut.mod_inv.mod_mul3/_122_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_157_ ));
 sky130_fd_sc_hd__xnor2_1 \uut.mod_inv.mod_mul3/_452_  (.A(\uut.mod_inv.mod_mul3/_156_ ),
    .B(\uut.mod_inv.mod_mul3/_157_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3/_158_ ));
 sky130_fd_sc_hd__xnor2_2 \uut.mod_inv.mod_mul3/_453_  (.A(\uut.mod_inv.mod_mul3/_048_ ),
    .B(\uut.mod_inv.mod_mul3/_158_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\uut.mod_inv.mod_mul3_out3[0] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.sh_mod1/_0_  (.A(\uut.mod_inv.sq_scl_in[0] ),
    .B(\uut.mod_inv.sq_scl_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out1[3] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.sh_mod1/_1_  (.A(\uut.mod_inv.sq_scl_in[1] ),
    .B(\uut.mod_inv.sq_scl_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out1[2] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.sh_mod1/_2_  (.A(\uut.mod_inv.sq_scl_in[0] ),
    .B(\uut.mod_inv.sq_scl_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out1[1] ));
 sky130_fd_sc_hd__clkbuf_1 \uut.mod_inv.sh_mod1/_3_  (.A(\uut.mod_inv.sq_scl_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out1[0] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.sh_mod2/_0_  (.A(\uut.mod_inv.sh1_xor_out[0] ),
    .B(\uut.mod_inv.sh1_xor_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out2[3] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.sh_mod2/_1_  (.A(\uut.mod_inv.sh1_xor_out[1] ),
    .B(\uut.mod_inv.sh1_xor_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out2[2] ));
 sky130_fd_sc_hd__xor2_1 \uut.mod_inv.sh_mod2/_2_  (.A(\uut.mod_inv.sh1_xor_out[0] ),
    .B(\uut.mod_inv.sh1_xor_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out2[1] ));
 sky130_fd_sc_hd__clkbuf_1 \uut.mod_inv.sh_mod2/_3_  (.A(\uut.mod_inv.sh1_xor_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uut.mod_inv.sq_scl_out2[0] ));
 assign uio_oe[0] = net36;
 assign uio_oe[1] = net37;
 assign uio_oe[2] = net38;
 assign uio_oe[3] = net39;
 assign uio_oe[4] = net40;
 assign uio_oe[5] = net41;
 assign uio_oe[6] = net42;
 assign uio_oe[7] = net43;
 assign uio_out[1] = net29;
 assign uio_out[2] = net30;
 assign uio_out[3] = net31;
 assign uio_out[4] = net32;
 assign uio_out[5] = net33;
 assign uio_out[6] = net34;
 assign uio_out[7] = net35;
endmodule
