VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_kianV_rv32ima_uLinux_SoC
  CLASS BLOCK ;
  FOREIGN tt_um_kianV_rv32ima_uLinux_SoC ;
  ORIGIN 0.000 0.000 ;
  SIZE 1359.760 BY 225.760 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.880 2.480 557.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.480 2.480 711.080 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.080 2.480 864.680 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1016.680 2.480 1018.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1170.280 2.480 1171.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.880 2.480 1325.480 223.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.680 2.480 634.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.280 2.480 787.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 939.880 2.480 941.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1093.480 2.480 1095.080 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1247.080 2.480 1248.680 223.280 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 145.670 224.760 145.970 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 148.430 224.760 148.730 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 142.910 224.760 143.210 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.390 224.760 137.690 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.630 224.760 134.930 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met4 ;
        RECT 131.870 224.760 132.170 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 126.350 224.760 126.650 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 123.590 224.760 123.890 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.830 224.760 121.130 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 115.310 224.760 115.610 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 112.550 224.760 112.850 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.790 224.760 110.090 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 104.270 224.760 104.570 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.510 224.760 101.810 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.750 224.760 99.050 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 49.070 224.760 49.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 46.310 224.760 46.610 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 43.550 224.760 43.850 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 38.030 224.760 38.330 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.270 224.760 35.570 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.510 224.760 32.810 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 71.150 224.760 71.450 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 68.390 224.760 68.690 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 65.630 224.760 65.930 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 60.110 224.760 60.410 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 57.350 224.760 57.650 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.590 224.760 54.890 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 93.230 224.760 93.530 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 90.470 224.760 90.770 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 87.710 224.760 88.010 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 82.190 224.760 82.490 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 79.430 224.760 79.730 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 76.670 224.760 76.970 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 221.625 1357.190 223.230 ;
        RECT 2.570 216.185 1357.190 219.015 ;
        RECT 2.570 210.745 1357.190 213.575 ;
        RECT 2.570 205.305 1357.190 208.135 ;
        RECT 2.570 199.865 1357.190 202.695 ;
        RECT 2.570 194.425 1357.190 197.255 ;
        RECT 2.570 188.985 1357.190 191.815 ;
        RECT 2.570 183.545 1357.190 186.375 ;
        RECT 2.570 178.105 1357.190 180.935 ;
        RECT 2.570 172.665 1357.190 175.495 ;
        RECT 2.570 167.225 1357.190 170.055 ;
        RECT 2.570 161.785 1357.190 164.615 ;
        RECT 2.570 156.345 1357.190 159.175 ;
        RECT 2.570 150.905 1357.190 153.735 ;
        RECT 2.570 145.465 1357.190 148.295 ;
        RECT 2.570 140.025 1357.190 142.855 ;
        RECT 2.570 134.585 1357.190 137.415 ;
        RECT 2.570 129.145 1357.190 131.975 ;
        RECT 2.570 123.705 1357.190 126.535 ;
        RECT 2.570 118.265 1357.190 121.095 ;
        RECT 2.570 112.825 1357.190 115.655 ;
        RECT 2.570 107.385 1357.190 110.215 ;
        RECT 2.570 101.945 1357.190 104.775 ;
        RECT 2.570 96.505 1357.190 99.335 ;
        RECT 2.570 91.065 1357.190 93.895 ;
        RECT 2.570 85.625 1357.190 88.455 ;
        RECT 2.570 80.185 1357.190 83.015 ;
        RECT 2.570 74.745 1357.190 77.575 ;
        RECT 2.570 69.305 1357.190 72.135 ;
        RECT 2.570 63.865 1357.190 66.695 ;
        RECT 2.570 58.425 1357.190 61.255 ;
        RECT 2.570 52.985 1357.190 55.815 ;
        RECT 2.570 47.545 1357.190 50.375 ;
        RECT 2.570 42.105 1357.190 44.935 ;
        RECT 2.570 36.665 1357.190 39.495 ;
        RECT 2.570 31.225 1357.190 34.055 ;
        RECT 2.570 25.785 1357.190 28.615 ;
        RECT 2.570 20.345 1357.190 23.175 ;
        RECT 2.570 14.905 1357.190 17.735 ;
        RECT 2.570 9.465 1357.190 12.295 ;
        RECT 2.570 4.025 1357.190 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 1357.000 223.125 ;
      LAYER met1 ;
        RECT 2.760 0.040 1357.000 225.720 ;
      LAYER met2 ;
        RECT 4.230 0.010 1354.140 225.750 ;
      LAYER met3 ;
        RECT 4.205 0.175 1350.035 225.585 ;
      LAYER met4 ;
        RECT 15.935 224.360 32.110 225.585 ;
        RECT 33.210 224.360 34.870 225.585 ;
        RECT 35.970 224.360 37.630 225.585 ;
        RECT 38.730 224.360 40.390 225.585 ;
        RECT 41.490 224.360 43.150 225.585 ;
        RECT 44.250 224.360 45.910 225.585 ;
        RECT 47.010 224.360 48.670 225.585 ;
        RECT 49.770 224.360 51.430 225.585 ;
        RECT 52.530 224.360 54.190 225.585 ;
        RECT 55.290 224.360 56.950 225.585 ;
        RECT 58.050 224.360 59.710 225.585 ;
        RECT 60.810 224.360 62.470 225.585 ;
        RECT 63.570 224.360 65.230 225.585 ;
        RECT 66.330 224.360 67.990 225.585 ;
        RECT 69.090 224.360 70.750 225.585 ;
        RECT 71.850 224.360 73.510 225.585 ;
        RECT 74.610 224.360 76.270 225.585 ;
        RECT 77.370 224.360 79.030 225.585 ;
        RECT 80.130 224.360 81.790 225.585 ;
        RECT 82.890 224.360 84.550 225.585 ;
        RECT 85.650 224.360 87.310 225.585 ;
        RECT 88.410 224.360 90.070 225.585 ;
        RECT 91.170 224.360 92.830 225.585 ;
        RECT 93.930 224.360 95.590 225.585 ;
        RECT 96.690 224.360 98.350 225.585 ;
        RECT 99.450 224.360 101.110 225.585 ;
        RECT 102.210 224.360 103.870 225.585 ;
        RECT 104.970 224.360 106.630 225.585 ;
        RECT 107.730 224.360 109.390 225.585 ;
        RECT 110.490 224.360 112.150 225.585 ;
        RECT 113.250 224.360 114.910 225.585 ;
        RECT 116.010 224.360 117.670 225.585 ;
        RECT 118.770 224.360 120.430 225.585 ;
        RECT 121.530 224.360 123.190 225.585 ;
        RECT 124.290 224.360 125.950 225.585 ;
        RECT 127.050 224.360 128.710 225.585 ;
        RECT 129.810 224.360 131.470 225.585 ;
        RECT 132.570 224.360 134.230 225.585 ;
        RECT 135.330 224.360 136.990 225.585 ;
        RECT 138.090 224.360 139.750 225.585 ;
        RECT 140.850 224.360 142.510 225.585 ;
        RECT 143.610 224.360 145.270 225.585 ;
        RECT 146.370 224.360 148.030 225.585 ;
        RECT 149.130 224.360 1306.105 225.585 ;
        RECT 15.935 223.680 1306.105 224.360 ;
        RECT 15.935 2.080 17.880 223.680 ;
        RECT 20.280 2.080 94.680 223.680 ;
        RECT 97.080 2.080 171.480 223.680 ;
        RECT 173.880 2.080 248.280 223.680 ;
        RECT 250.680 2.080 325.080 223.680 ;
        RECT 327.480 2.080 401.880 223.680 ;
        RECT 404.280 2.080 478.680 223.680 ;
        RECT 481.080 2.080 555.480 223.680 ;
        RECT 557.880 2.080 632.280 223.680 ;
        RECT 634.680 2.080 709.080 223.680 ;
        RECT 711.480 2.080 785.880 223.680 ;
        RECT 788.280 2.080 862.680 223.680 ;
        RECT 865.080 2.080 939.480 223.680 ;
        RECT 941.880 2.080 1016.280 223.680 ;
        RECT 1018.680 2.080 1093.080 223.680 ;
        RECT 1095.480 2.080 1169.880 223.680 ;
        RECT 1172.280 2.080 1246.680 223.680 ;
        RECT 1249.080 2.080 1306.105 223.680 ;
        RECT 15.935 0.855 1306.105 2.080 ;
  END
END tt_um_kianV_rv32ima_uLinux_SoC
END LIBRARY

