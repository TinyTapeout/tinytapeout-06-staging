VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_analog_test
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_analog_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 0.000 2.500 225.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 0.000 50.500 225.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 95.970 24.030 96.300 24.200 ;
        RECT 96.510 24.030 96.840 24.200 ;
        RECT 97.050 24.030 97.380 24.200 ;
        RECT 97.590 24.030 97.920 24.200 ;
        RECT 98.130 24.030 98.460 24.200 ;
        RECT 96.050 22.215 96.220 24.030 ;
        RECT 96.590 22.215 96.760 24.030 ;
        RECT 97.130 22.215 97.300 24.030 ;
        RECT 97.670 22.215 97.840 24.030 ;
        RECT 98.210 22.215 98.380 24.030 ;
        RECT 96.050 18.580 96.220 20.395 ;
        RECT 96.590 18.580 96.760 20.395 ;
        RECT 97.130 18.580 97.300 20.395 ;
        RECT 97.670 18.580 97.840 20.395 ;
        RECT 98.210 18.580 98.380 20.395 ;
        RECT 95.970 18.410 96.300 18.580 ;
        RECT 96.510 18.410 96.840 18.580 ;
        RECT 97.050 18.410 97.380 18.580 ;
        RECT 97.590 18.410 97.920 18.580 ;
        RECT 98.130 18.410 98.460 18.580 ;
      LAYER mcon ;
        RECT 96.050 18.410 96.220 20.395 ;
        RECT 96.590 18.410 96.760 20.395 ;
        RECT 97.130 18.410 97.300 20.395 ;
        RECT 97.670 18.410 97.840 20.395 ;
        RECT 98.210 18.410 98.380 20.395 ;
      LAYER met1 ;
        RECT 94.000 26.570 96.160 33.020 ;
        RECT 94.990 25.980 95.290 26.570 ;
        RECT 94.990 25.680 96.310 25.980 ;
        RECT 96.010 24.280 96.310 25.680 ;
        RECT 95.970 24.200 96.310 24.280 ;
        RECT 96.560 24.200 96.790 24.260 ;
        RECT 97.100 24.200 97.330 24.260 ;
        RECT 97.640 24.200 97.870 24.260 ;
        RECT 98.180 24.200 98.410 24.260 ;
        RECT 95.920 22.580 98.560 24.200 ;
        RECT 96.020 22.155 96.250 22.580 ;
        RECT 96.560 22.155 96.790 22.580 ;
        RECT 97.100 22.155 97.330 22.580 ;
        RECT 97.640 22.155 97.870 22.580 ;
        RECT 98.180 22.155 98.410 22.580 ;
        RECT 96.020 19.850 96.250 20.455 ;
        RECT 96.560 19.850 96.790 20.455 ;
        RECT 95.930 8.365 96.880 19.850 ;
        RECT 97.100 19.820 97.330 20.455 ;
        RECT 97.640 19.820 97.870 20.455 ;
        RECT 98.180 19.820 98.410 20.455 ;
        RECT 97.050 13.520 98.450 19.820 ;
        RECT 97.050 12.120 155.700 13.520 ;
        RECT 123.570 8.365 125.980 8.650 ;
        RECT 154.300 8.380 155.700 12.120 ;
        RECT 95.930 7.415 125.980 8.365 ;
        RECT 123.570 6.610 125.980 7.415 ;
        RECT 154.130 6.830 155.910 8.380 ;
        RECT 154.300 6.300 155.700 6.830 ;
      LAYER via ;
        RECT 94.150 30.950 95.950 32.600 ;
        RECT 123.620 6.610 125.930 8.650 ;
        RECT 154.180 6.830 155.860 8.380 ;
      LAYER met2 ;
        RECT 94.150 30.900 95.950 32.650 ;
        RECT 123.620 6.560 125.930 8.700 ;
        RECT 154.180 6.780 155.860 8.430 ;
      LAYER via2 ;
        RECT 94.150 30.950 95.950 32.600 ;
        RECT 123.620 6.610 125.930 8.650 ;
        RECT 154.180 6.830 155.860 8.380 ;
      LAYER met3 ;
        RECT 94.100 30.925 96.000 32.625 ;
        RECT 123.570 6.585 125.980 8.675 ;
        RECT 154.130 6.805 155.910 8.405 ;
      LAYER via3 ;
        RECT 94.150 30.950 95.950 32.600 ;
        RECT 123.620 6.610 125.930 8.650 ;
        RECT 154.180 6.830 155.860 8.380 ;
      LAYER met4 ;
        RECT 48.810 30.780 49.000 32.850 ;
        RECT 50.500 30.780 96.300 32.850 ;
        RECT 123.615 6.605 125.935 8.655 ;
        RECT 154.175 6.825 155.865 8.385 ;
        RECT 124.540 6.220 125.140 6.605 ;
        RECT 124.540 5.620 135.080 6.220 ;
        RECT 134.480 1.000 135.080 5.620 ;
        RECT 154.690 4.100 155.290 6.825 ;
        RECT 154.690 3.500 157.160 4.100 ;
        RECT 156.560 1.000 157.160 3.500 ;
  END
END tt_um_mattvenn_analog_test
END LIBRARY

