module tt_um_gfg_development_tros_dup (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire data_stream;
 wire \ena_syncs[0] ;
 wire \ena_syncs[1] ;
 wire \ena_syncs[2] ;
 wire \fmeasurment_einv_sub_ros.counts[0] ;
 wire \fmeasurment_einv_sub_ros.counts[10] ;
 wire \fmeasurment_einv_sub_ros.counts[11] ;
 wire \fmeasurment_einv_sub_ros.counts[12] ;
 wire \fmeasurment_einv_sub_ros.counts[13] ;
 wire \fmeasurment_einv_sub_ros.counts[14] ;
 wire \fmeasurment_einv_sub_ros.counts[15] ;
 wire \fmeasurment_einv_sub_ros.counts[16] ;
 wire \fmeasurment_einv_sub_ros.counts[17] ;
 wire \fmeasurment_einv_sub_ros.counts[18] ;
 wire \fmeasurment_einv_sub_ros.counts[19] ;
 wire \fmeasurment_einv_sub_ros.counts[1] ;
 wire \fmeasurment_einv_sub_ros.counts[2] ;
 wire \fmeasurment_einv_sub_ros.counts[3] ;
 wire \fmeasurment_einv_sub_ros.counts[4] ;
 wire \fmeasurment_einv_sub_ros.counts[5] ;
 wire \fmeasurment_einv_sub_ros.counts[6] ;
 wire \fmeasurment_einv_sub_ros.counts[7] ;
 wire \fmeasurment_einv_sub_ros.counts[8] ;
 wire \fmeasurment_einv_sub_ros.counts[9] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[0] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[10] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[11] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[12] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[13] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[14] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[15] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[16] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[17] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[18] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[19] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[1] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[2] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[3] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[4] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[5] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[6] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[7] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[8] ;
 wire \fmeasurment_einv_sub_ros.cycle_count[9] ;
 wire \fmeasurment_einv_sub_ros.divided_clk ;
 wire \fmeasurment_einv_sub_ros.latch_counter_syncs[0] ;
 wire \fmeasurment_einv_sub_ros.latch_counter_syncs[1] ;
 wire \fmeasurment_einv_sub_ros.latch_counter_syncs[2] ;
 wire \fmeasurment_einv_sub_ros.reset_syncs[0] ;
 wire \fmeasurment_einv_sub_ros.reset_syncs[1] ;
 wire \fmeasurment_einv_sub_ros.reset_syncs[2] ;
 wire \fmeasurment_nand4_cap_ros.counts[0] ;
 wire \fmeasurment_nand4_cap_ros.counts[10] ;
 wire \fmeasurment_nand4_cap_ros.counts[11] ;
 wire \fmeasurment_nand4_cap_ros.counts[12] ;
 wire \fmeasurment_nand4_cap_ros.counts[13] ;
 wire \fmeasurment_nand4_cap_ros.counts[14] ;
 wire \fmeasurment_nand4_cap_ros.counts[15] ;
 wire \fmeasurment_nand4_cap_ros.counts[16] ;
 wire \fmeasurment_nand4_cap_ros.counts[17] ;
 wire \fmeasurment_nand4_cap_ros.counts[18] ;
 wire \fmeasurment_nand4_cap_ros.counts[19] ;
 wire \fmeasurment_nand4_cap_ros.counts[1] ;
 wire \fmeasurment_nand4_cap_ros.counts[2] ;
 wire \fmeasurment_nand4_cap_ros.counts[3] ;
 wire \fmeasurment_nand4_cap_ros.counts[4] ;
 wire \fmeasurment_nand4_cap_ros.counts[5] ;
 wire \fmeasurment_nand4_cap_ros.counts[6] ;
 wire \fmeasurment_nand4_cap_ros.counts[7] ;
 wire \fmeasurment_nand4_cap_ros.counts[8] ;
 wire \fmeasurment_nand4_cap_ros.counts[9] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[0] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[10] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[11] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[12] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[13] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[14] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[15] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[16] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[17] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[18] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[19] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[1] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[2] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[3] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[4] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[5] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[6] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[7] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[8] ;
 wire \fmeasurment_nand4_cap_ros.cycle_count[9] ;
 wire \fmeasurment_nand4_cap_ros.divided_clk ;
 wire \fmeasurment_nand4_cap_ros.latch_counter_syncs[0] ;
 wire \fmeasurment_nand4_cap_ros.latch_counter_syncs[1] ;
 wire \fmeasurment_nand4_cap_ros.latch_counter_syncs[2] ;
 wire \fmeasurment_nand4_cap_ros.reset_syncs[0] ;
 wire \fmeasurment_nand4_cap_ros.reset_syncs[1] ;
 wire \fmeasurment_nand4_cap_ros.reset_syncs[2] ;
 wire \fmeasurment_nand4_ros.counts[0] ;
 wire \fmeasurment_nand4_ros.counts[10] ;
 wire \fmeasurment_nand4_ros.counts[11] ;
 wire \fmeasurment_nand4_ros.counts[12] ;
 wire \fmeasurment_nand4_ros.counts[13] ;
 wire \fmeasurment_nand4_ros.counts[14] ;
 wire \fmeasurment_nand4_ros.counts[15] ;
 wire \fmeasurment_nand4_ros.counts[16] ;
 wire \fmeasurment_nand4_ros.counts[17] ;
 wire \fmeasurment_nand4_ros.counts[18] ;
 wire \fmeasurment_nand4_ros.counts[19] ;
 wire \fmeasurment_nand4_ros.counts[1] ;
 wire \fmeasurment_nand4_ros.counts[2] ;
 wire \fmeasurment_nand4_ros.counts[3] ;
 wire \fmeasurment_nand4_ros.counts[4] ;
 wire \fmeasurment_nand4_ros.counts[5] ;
 wire \fmeasurment_nand4_ros.counts[6] ;
 wire \fmeasurment_nand4_ros.counts[7] ;
 wire \fmeasurment_nand4_ros.counts[8] ;
 wire \fmeasurment_nand4_ros.counts[9] ;
 wire \fmeasurment_nand4_ros.cycle_count[0] ;
 wire \fmeasurment_nand4_ros.cycle_count[10] ;
 wire \fmeasurment_nand4_ros.cycle_count[11] ;
 wire \fmeasurment_nand4_ros.cycle_count[12] ;
 wire \fmeasurment_nand4_ros.cycle_count[13] ;
 wire \fmeasurment_nand4_ros.cycle_count[14] ;
 wire \fmeasurment_nand4_ros.cycle_count[15] ;
 wire \fmeasurment_nand4_ros.cycle_count[16] ;
 wire \fmeasurment_nand4_ros.cycle_count[17] ;
 wire \fmeasurment_nand4_ros.cycle_count[18] ;
 wire \fmeasurment_nand4_ros.cycle_count[19] ;
 wire \fmeasurment_nand4_ros.cycle_count[1] ;
 wire \fmeasurment_nand4_ros.cycle_count[2] ;
 wire \fmeasurment_nand4_ros.cycle_count[3] ;
 wire \fmeasurment_nand4_ros.cycle_count[4] ;
 wire \fmeasurment_nand4_ros.cycle_count[5] ;
 wire \fmeasurment_nand4_ros.cycle_count[6] ;
 wire \fmeasurment_nand4_ros.cycle_count[7] ;
 wire \fmeasurment_nand4_ros.cycle_count[8] ;
 wire \fmeasurment_nand4_ros.cycle_count[9] ;
 wire \fmeasurment_nand4_ros.divided_clk ;
 wire \fmeasurment_nand4_ros.latch_counter_syncs[0] ;
 wire \fmeasurment_nand4_ros.latch_counter_syncs[1] ;
 wire \fmeasurment_nand4_ros.latch_counter_syncs[2] ;
 wire \fmeasurment_nand4_ros.reset_syncs[0] ;
 wire \fmeasurment_nand4_ros.reset_syncs[1] ;
 wire \fmeasurment_nand4_ros.reset_syncs[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \ros_einv_sub.nets_notouch_[0] ;
 wire \ros_einv_sub.nets_notouch_[10] ;
 wire \ros_einv_sub.nets_notouch_[11] ;
 wire \ros_einv_sub.nets_notouch_[12] ;
 wire \ros_einv_sub.nets_notouch_[13] ;
 wire \ros_einv_sub.nets_notouch_[14] ;
 wire \ros_einv_sub.nets_notouch_[15] ;
 wire \ros_einv_sub.nets_notouch_[16] ;
 wire \ros_einv_sub.nets_notouch_[17] ;
 wire \ros_einv_sub.nets_notouch_[18] ;
 wire \ros_einv_sub.nets_notouch_[19] ;
 wire \ros_einv_sub.nets_notouch_[1] ;
 wire \ros_einv_sub.nets_notouch_[20] ;
 wire \ros_einv_sub.nets_notouch_[21] ;
 wire \ros_einv_sub.nets_notouch_[22] ;
 wire \ros_einv_sub.nets_notouch_[23] ;
 wire \ros_einv_sub.nets_notouch_[24] ;
 wire \ros_einv_sub.nets_notouch_[2] ;
 wire \ros_einv_sub.nets_notouch_[3] ;
 wire \ros_einv_sub.nets_notouch_[4] ;
 wire \ros_einv_sub.nets_notouch_[5] ;
 wire \ros_einv_sub.nets_notouch_[6] ;
 wire \ros_einv_sub.nets_notouch_[7] ;
 wire \ros_einv_sub.nets_notouch_[8] ;
 wire \ros_einv_sub.nets_notouch_[9] ;
 wire \ros_einv_sub.sub_voltage_notouch_ ;
 wire \ros_nand4.nets_notouch_[0] ;
 wire \ros_nand4.nets_notouch_[10] ;
 wire \ros_nand4.nets_notouch_[11] ;
 wire \ros_nand4.nets_notouch_[12] ;
 wire \ros_nand4.nets_notouch_[13] ;
 wire \ros_nand4.nets_notouch_[14] ;
 wire \ros_nand4.nets_notouch_[15] ;
 wire \ros_nand4.nets_notouch_[16] ;
 wire \ros_nand4.nets_notouch_[17] ;
 wire \ros_nand4.nets_notouch_[18] ;
 wire \ros_nand4.nets_notouch_[19] ;
 wire \ros_nand4.nets_notouch_[1] ;
 wire \ros_nand4.nets_notouch_[20] ;
 wire \ros_nand4.nets_notouch_[21] ;
 wire \ros_nand4.nets_notouch_[22] ;
 wire \ros_nand4.nets_notouch_[23] ;
 wire \ros_nand4.nets_notouch_[24] ;
 wire \ros_nand4.nets_notouch_[25] ;
 wire \ros_nand4.nets_notouch_[26] ;
 wire \ros_nand4.nets_notouch_[27] ;
 wire \ros_nand4.nets_notouch_[28] ;
 wire \ros_nand4.nets_notouch_[29] ;
 wire \ros_nand4.nets_notouch_[2] ;
 wire \ros_nand4.nets_notouch_[30] ;
 wire \ros_nand4.nets_notouch_[31] ;
 wire \ros_nand4.nets_notouch_[32] ;
 wire \ros_nand4.nets_notouch_[33] ;
 wire \ros_nand4.nets_notouch_[34] ;
 wire \ros_nand4.nets_notouch_[35] ;
 wire \ros_nand4.nets_notouch_[36] ;
 wire \ros_nand4.nets_notouch_[37] ;
 wire \ros_nand4.nets_notouch_[38] ;
 wire \ros_nand4.nets_notouch_[39] ;
 wire \ros_nand4.nets_notouch_[3] ;
 wire \ros_nand4.nets_notouch_[40] ;
 wire \ros_nand4.nets_notouch_[41] ;
 wire \ros_nand4.nets_notouch_[42] ;
 wire \ros_nand4.nets_notouch_[43] ;
 wire \ros_nand4.nets_notouch_[44] ;
 wire \ros_nand4.nets_notouch_[45] ;
 wire \ros_nand4.nets_notouch_[46] ;
 wire \ros_nand4.nets_notouch_[47] ;
 wire \ros_nand4.nets_notouch_[48] ;
 wire \ros_nand4.nets_notouch_[49] ;
 wire \ros_nand4.nets_notouch_[4] ;
 wire \ros_nand4.nets_notouch_[50] ;
 wire \ros_nand4.nets_notouch_[51] ;
 wire \ros_nand4.nets_notouch_[52] ;
 wire \ros_nand4.nets_notouch_[53] ;
 wire \ros_nand4.nets_notouch_[54] ;
 wire \ros_nand4.nets_notouch_[55] ;
 wire \ros_nand4.nets_notouch_[56] ;
 wire \ros_nand4.nets_notouch_[57] ;
 wire \ros_nand4.nets_notouch_[58] ;
 wire \ros_nand4.nets_notouch_[59] ;
 wire \ros_nand4.nets_notouch_[5] ;
 wire \ros_nand4.nets_notouch_[60] ;
 wire \ros_nand4.nets_notouch_[61] ;
 wire \ros_nand4.nets_notouch_[62] ;
 wire \ros_nand4.nets_notouch_[63] ;
 wire \ros_nand4.nets_notouch_[64] ;
 wire \ros_nand4.nets_notouch_[65] ;
 wire \ros_nand4.nets_notouch_[66] ;
 wire \ros_nand4.nets_notouch_[6] ;
 wire \ros_nand4.nets_notouch_[7] ;
 wire \ros_nand4.nets_notouch_[8] ;
 wire \ros_nand4.nets_notouch_[9] ;
 wire \ros_nand4_cap.nets_notouch_[0] ;
 wire \ros_nand4_cap.nets_notouch_[10] ;
 wire \ros_nand4_cap.nets_notouch_[11] ;
 wire \ros_nand4_cap.nets_notouch_[12] ;
 wire \ros_nand4_cap.nets_notouch_[13] ;
 wire \ros_nand4_cap.nets_notouch_[14] ;
 wire \ros_nand4_cap.nets_notouch_[15] ;
 wire \ros_nand4_cap.nets_notouch_[16] ;
 wire \ros_nand4_cap.nets_notouch_[17] ;
 wire \ros_nand4_cap.nets_notouch_[18] ;
 wire \ros_nand4_cap.nets_notouch_[19] ;
 wire \ros_nand4_cap.nets_notouch_[1] ;
 wire \ros_nand4_cap.nets_notouch_[20] ;
 wire \ros_nand4_cap.nets_notouch_[21] ;
 wire \ros_nand4_cap.nets_notouch_[22] ;
 wire \ros_nand4_cap.nets_notouch_[23] ;
 wire \ros_nand4_cap.nets_notouch_[24] ;
 wire \ros_nand4_cap.nets_notouch_[25] ;
 wire \ros_nand4_cap.nets_notouch_[26] ;
 wire \ros_nand4_cap.nets_notouch_[27] ;
 wire \ros_nand4_cap.nets_notouch_[28] ;
 wire \ros_nand4_cap.nets_notouch_[29] ;
 wire \ros_nand4_cap.nets_notouch_[2] ;
 wire \ros_nand4_cap.nets_notouch_[30] ;
 wire \ros_nand4_cap.nets_notouch_[31] ;
 wire \ros_nand4_cap.nets_notouch_[32] ;
 wire \ros_nand4_cap.nets_notouch_[33] ;
 wire \ros_nand4_cap.nets_notouch_[34] ;
 wire \ros_nand4_cap.nets_notouch_[3] ;
 wire \ros_nand4_cap.nets_notouch_[4] ;
 wire \ros_nand4_cap.nets_notouch_[5] ;
 wire \ros_nand4_cap.nets_notouch_[6] ;
 wire \ros_nand4_cap.nets_notouch_[7] ;
 wire \ros_nand4_cap.nets_notouch_[8] ;
 wire \ros_nand4_cap.nets_notouch_[9] ;
 wire \ros_nand4_cap.open_nets_notouch_[0] ;
 wire \ros_nand4_cap.open_nets_notouch_[100] ;
 wire \ros_nand4_cap.open_nets_notouch_[101] ;
 wire \ros_nand4_cap.open_nets_notouch_[102] ;
 wire \ros_nand4_cap.open_nets_notouch_[103] ;
 wire \ros_nand4_cap.open_nets_notouch_[104] ;
 wire \ros_nand4_cap.open_nets_notouch_[105] ;
 wire \ros_nand4_cap.open_nets_notouch_[106] ;
 wire \ros_nand4_cap.open_nets_notouch_[107] ;
 wire \ros_nand4_cap.open_nets_notouch_[108] ;
 wire \ros_nand4_cap.open_nets_notouch_[109] ;
 wire \ros_nand4_cap.open_nets_notouch_[10] ;
 wire \ros_nand4_cap.open_nets_notouch_[110] ;
 wire \ros_nand4_cap.open_nets_notouch_[111] ;
 wire \ros_nand4_cap.open_nets_notouch_[112] ;
 wire \ros_nand4_cap.open_nets_notouch_[113] ;
 wire \ros_nand4_cap.open_nets_notouch_[114] ;
 wire \ros_nand4_cap.open_nets_notouch_[115] ;
 wire \ros_nand4_cap.open_nets_notouch_[116] ;
 wire \ros_nand4_cap.open_nets_notouch_[117] ;
 wire \ros_nand4_cap.open_nets_notouch_[118] ;
 wire \ros_nand4_cap.open_nets_notouch_[119] ;
 wire \ros_nand4_cap.open_nets_notouch_[11] ;
 wire \ros_nand4_cap.open_nets_notouch_[120] ;
 wire \ros_nand4_cap.open_nets_notouch_[121] ;
 wire \ros_nand4_cap.open_nets_notouch_[122] ;
 wire \ros_nand4_cap.open_nets_notouch_[123] ;
 wire \ros_nand4_cap.open_nets_notouch_[124] ;
 wire \ros_nand4_cap.open_nets_notouch_[125] ;
 wire \ros_nand4_cap.open_nets_notouch_[126] ;
 wire \ros_nand4_cap.open_nets_notouch_[127] ;
 wire \ros_nand4_cap.open_nets_notouch_[128] ;
 wire \ros_nand4_cap.open_nets_notouch_[129] ;
 wire \ros_nand4_cap.open_nets_notouch_[12] ;
 wire \ros_nand4_cap.open_nets_notouch_[130] ;
 wire \ros_nand4_cap.open_nets_notouch_[131] ;
 wire \ros_nand4_cap.open_nets_notouch_[132] ;
 wire \ros_nand4_cap.open_nets_notouch_[133] ;
 wire \ros_nand4_cap.open_nets_notouch_[134] ;
 wire \ros_nand4_cap.open_nets_notouch_[135] ;
 wire \ros_nand4_cap.open_nets_notouch_[136] ;
 wire \ros_nand4_cap.open_nets_notouch_[137] ;
 wire \ros_nand4_cap.open_nets_notouch_[138] ;
 wire \ros_nand4_cap.open_nets_notouch_[139] ;
 wire \ros_nand4_cap.open_nets_notouch_[13] ;
 wire \ros_nand4_cap.open_nets_notouch_[140] ;
 wire \ros_nand4_cap.open_nets_notouch_[141] ;
 wire \ros_nand4_cap.open_nets_notouch_[142] ;
 wire \ros_nand4_cap.open_nets_notouch_[143] ;
 wire \ros_nand4_cap.open_nets_notouch_[144] ;
 wire \ros_nand4_cap.open_nets_notouch_[145] ;
 wire \ros_nand4_cap.open_nets_notouch_[146] ;
 wire \ros_nand4_cap.open_nets_notouch_[147] ;
 wire \ros_nand4_cap.open_nets_notouch_[148] ;
 wire \ros_nand4_cap.open_nets_notouch_[149] ;
 wire \ros_nand4_cap.open_nets_notouch_[14] ;
 wire \ros_nand4_cap.open_nets_notouch_[150] ;
 wire \ros_nand4_cap.open_nets_notouch_[151] ;
 wire \ros_nand4_cap.open_nets_notouch_[152] ;
 wire \ros_nand4_cap.open_nets_notouch_[153] ;
 wire \ros_nand4_cap.open_nets_notouch_[154] ;
 wire \ros_nand4_cap.open_nets_notouch_[155] ;
 wire \ros_nand4_cap.open_nets_notouch_[156] ;
 wire \ros_nand4_cap.open_nets_notouch_[157] ;
 wire \ros_nand4_cap.open_nets_notouch_[158] ;
 wire \ros_nand4_cap.open_nets_notouch_[159] ;
 wire \ros_nand4_cap.open_nets_notouch_[15] ;
 wire \ros_nand4_cap.open_nets_notouch_[160] ;
 wire \ros_nand4_cap.open_nets_notouch_[161] ;
 wire \ros_nand4_cap.open_nets_notouch_[162] ;
 wire \ros_nand4_cap.open_nets_notouch_[163] ;
 wire \ros_nand4_cap.open_nets_notouch_[164] ;
 wire \ros_nand4_cap.open_nets_notouch_[165] ;
 wire \ros_nand4_cap.open_nets_notouch_[166] ;
 wire \ros_nand4_cap.open_nets_notouch_[167] ;
 wire \ros_nand4_cap.open_nets_notouch_[168] ;
 wire \ros_nand4_cap.open_nets_notouch_[169] ;
 wire \ros_nand4_cap.open_nets_notouch_[16] ;
 wire \ros_nand4_cap.open_nets_notouch_[170] ;
 wire \ros_nand4_cap.open_nets_notouch_[171] ;
 wire \ros_nand4_cap.open_nets_notouch_[172] ;
 wire \ros_nand4_cap.open_nets_notouch_[173] ;
 wire \ros_nand4_cap.open_nets_notouch_[174] ;
 wire \ros_nand4_cap.open_nets_notouch_[175] ;
 wire \ros_nand4_cap.open_nets_notouch_[176] ;
 wire \ros_nand4_cap.open_nets_notouch_[177] ;
 wire \ros_nand4_cap.open_nets_notouch_[178] ;
 wire \ros_nand4_cap.open_nets_notouch_[179] ;
 wire \ros_nand4_cap.open_nets_notouch_[17] ;
 wire \ros_nand4_cap.open_nets_notouch_[180] ;
 wire \ros_nand4_cap.open_nets_notouch_[181] ;
 wire \ros_nand4_cap.open_nets_notouch_[182] ;
 wire \ros_nand4_cap.open_nets_notouch_[183] ;
 wire \ros_nand4_cap.open_nets_notouch_[184] ;
 wire \ros_nand4_cap.open_nets_notouch_[185] ;
 wire \ros_nand4_cap.open_nets_notouch_[186] ;
 wire \ros_nand4_cap.open_nets_notouch_[187] ;
 wire \ros_nand4_cap.open_nets_notouch_[188] ;
 wire \ros_nand4_cap.open_nets_notouch_[189] ;
 wire \ros_nand4_cap.open_nets_notouch_[18] ;
 wire \ros_nand4_cap.open_nets_notouch_[190] ;
 wire \ros_nand4_cap.open_nets_notouch_[191] ;
 wire \ros_nand4_cap.open_nets_notouch_[192] ;
 wire \ros_nand4_cap.open_nets_notouch_[193] ;
 wire \ros_nand4_cap.open_nets_notouch_[194] ;
 wire \ros_nand4_cap.open_nets_notouch_[195] ;
 wire \ros_nand4_cap.open_nets_notouch_[196] ;
 wire \ros_nand4_cap.open_nets_notouch_[197] ;
 wire \ros_nand4_cap.open_nets_notouch_[198] ;
 wire \ros_nand4_cap.open_nets_notouch_[199] ;
 wire \ros_nand4_cap.open_nets_notouch_[19] ;
 wire \ros_nand4_cap.open_nets_notouch_[1] ;
 wire \ros_nand4_cap.open_nets_notouch_[200] ;
 wire \ros_nand4_cap.open_nets_notouch_[201] ;
 wire \ros_nand4_cap.open_nets_notouch_[202] ;
 wire \ros_nand4_cap.open_nets_notouch_[203] ;
 wire \ros_nand4_cap.open_nets_notouch_[204] ;
 wire \ros_nand4_cap.open_nets_notouch_[205] ;
 wire \ros_nand4_cap.open_nets_notouch_[206] ;
 wire \ros_nand4_cap.open_nets_notouch_[207] ;
 wire \ros_nand4_cap.open_nets_notouch_[208] ;
 wire \ros_nand4_cap.open_nets_notouch_[209] ;
 wire \ros_nand4_cap.open_nets_notouch_[20] ;
 wire \ros_nand4_cap.open_nets_notouch_[210] ;
 wire \ros_nand4_cap.open_nets_notouch_[211] ;
 wire \ros_nand4_cap.open_nets_notouch_[212] ;
 wire \ros_nand4_cap.open_nets_notouch_[213] ;
 wire \ros_nand4_cap.open_nets_notouch_[214] ;
 wire \ros_nand4_cap.open_nets_notouch_[215] ;
 wire \ros_nand4_cap.open_nets_notouch_[216] ;
 wire \ros_nand4_cap.open_nets_notouch_[217] ;
 wire \ros_nand4_cap.open_nets_notouch_[218] ;
 wire \ros_nand4_cap.open_nets_notouch_[219] ;
 wire \ros_nand4_cap.open_nets_notouch_[21] ;
 wire \ros_nand4_cap.open_nets_notouch_[220] ;
 wire \ros_nand4_cap.open_nets_notouch_[221] ;
 wire \ros_nand4_cap.open_nets_notouch_[222] ;
 wire \ros_nand4_cap.open_nets_notouch_[223] ;
 wire \ros_nand4_cap.open_nets_notouch_[224] ;
 wire \ros_nand4_cap.open_nets_notouch_[225] ;
 wire \ros_nand4_cap.open_nets_notouch_[226] ;
 wire \ros_nand4_cap.open_nets_notouch_[227] ;
 wire \ros_nand4_cap.open_nets_notouch_[228] ;
 wire \ros_nand4_cap.open_nets_notouch_[229] ;
 wire \ros_nand4_cap.open_nets_notouch_[22] ;
 wire \ros_nand4_cap.open_nets_notouch_[230] ;
 wire \ros_nand4_cap.open_nets_notouch_[231] ;
 wire \ros_nand4_cap.open_nets_notouch_[232] ;
 wire \ros_nand4_cap.open_nets_notouch_[233] ;
 wire \ros_nand4_cap.open_nets_notouch_[234] ;
 wire \ros_nand4_cap.open_nets_notouch_[235] ;
 wire \ros_nand4_cap.open_nets_notouch_[236] ;
 wire \ros_nand4_cap.open_nets_notouch_[237] ;
 wire \ros_nand4_cap.open_nets_notouch_[238] ;
 wire \ros_nand4_cap.open_nets_notouch_[239] ;
 wire \ros_nand4_cap.open_nets_notouch_[23] ;
 wire \ros_nand4_cap.open_nets_notouch_[240] ;
 wire \ros_nand4_cap.open_nets_notouch_[241] ;
 wire \ros_nand4_cap.open_nets_notouch_[242] ;
 wire \ros_nand4_cap.open_nets_notouch_[243] ;
 wire \ros_nand4_cap.open_nets_notouch_[244] ;
 wire \ros_nand4_cap.open_nets_notouch_[245] ;
 wire \ros_nand4_cap.open_nets_notouch_[246] ;
 wire \ros_nand4_cap.open_nets_notouch_[247] ;
 wire \ros_nand4_cap.open_nets_notouch_[248] ;
 wire \ros_nand4_cap.open_nets_notouch_[249] ;
 wire \ros_nand4_cap.open_nets_notouch_[24] ;
 wire \ros_nand4_cap.open_nets_notouch_[250] ;
 wire \ros_nand4_cap.open_nets_notouch_[251] ;
 wire \ros_nand4_cap.open_nets_notouch_[252] ;
 wire \ros_nand4_cap.open_nets_notouch_[253] ;
 wire \ros_nand4_cap.open_nets_notouch_[254] ;
 wire \ros_nand4_cap.open_nets_notouch_[255] ;
 wire \ros_nand4_cap.open_nets_notouch_[256] ;
 wire \ros_nand4_cap.open_nets_notouch_[257] ;
 wire \ros_nand4_cap.open_nets_notouch_[258] ;
 wire \ros_nand4_cap.open_nets_notouch_[259] ;
 wire \ros_nand4_cap.open_nets_notouch_[25] ;
 wire \ros_nand4_cap.open_nets_notouch_[260] ;
 wire \ros_nand4_cap.open_nets_notouch_[261] ;
 wire \ros_nand4_cap.open_nets_notouch_[262] ;
 wire \ros_nand4_cap.open_nets_notouch_[263] ;
 wire \ros_nand4_cap.open_nets_notouch_[264] ;
 wire \ros_nand4_cap.open_nets_notouch_[265] ;
 wire \ros_nand4_cap.open_nets_notouch_[266] ;
 wire \ros_nand4_cap.open_nets_notouch_[267] ;
 wire \ros_nand4_cap.open_nets_notouch_[268] ;
 wire \ros_nand4_cap.open_nets_notouch_[269] ;
 wire \ros_nand4_cap.open_nets_notouch_[26] ;
 wire \ros_nand4_cap.open_nets_notouch_[270] ;
 wire \ros_nand4_cap.open_nets_notouch_[271] ;
 wire \ros_nand4_cap.open_nets_notouch_[272] ;
 wire \ros_nand4_cap.open_nets_notouch_[273] ;
 wire \ros_nand4_cap.open_nets_notouch_[274] ;
 wire \ros_nand4_cap.open_nets_notouch_[275] ;
 wire \ros_nand4_cap.open_nets_notouch_[276] ;
 wire \ros_nand4_cap.open_nets_notouch_[277] ;
 wire \ros_nand4_cap.open_nets_notouch_[278] ;
 wire \ros_nand4_cap.open_nets_notouch_[279] ;
 wire \ros_nand4_cap.open_nets_notouch_[27] ;
 wire \ros_nand4_cap.open_nets_notouch_[28] ;
 wire \ros_nand4_cap.open_nets_notouch_[29] ;
 wire \ros_nand4_cap.open_nets_notouch_[2] ;
 wire \ros_nand4_cap.open_nets_notouch_[30] ;
 wire \ros_nand4_cap.open_nets_notouch_[31] ;
 wire \ros_nand4_cap.open_nets_notouch_[32] ;
 wire \ros_nand4_cap.open_nets_notouch_[33] ;
 wire \ros_nand4_cap.open_nets_notouch_[34] ;
 wire \ros_nand4_cap.open_nets_notouch_[35] ;
 wire \ros_nand4_cap.open_nets_notouch_[36] ;
 wire \ros_nand4_cap.open_nets_notouch_[37] ;
 wire \ros_nand4_cap.open_nets_notouch_[38] ;
 wire \ros_nand4_cap.open_nets_notouch_[39] ;
 wire \ros_nand4_cap.open_nets_notouch_[3] ;
 wire \ros_nand4_cap.open_nets_notouch_[40] ;
 wire \ros_nand4_cap.open_nets_notouch_[41] ;
 wire \ros_nand4_cap.open_nets_notouch_[42] ;
 wire \ros_nand4_cap.open_nets_notouch_[43] ;
 wire \ros_nand4_cap.open_nets_notouch_[44] ;
 wire \ros_nand4_cap.open_nets_notouch_[45] ;
 wire \ros_nand4_cap.open_nets_notouch_[46] ;
 wire \ros_nand4_cap.open_nets_notouch_[47] ;
 wire \ros_nand4_cap.open_nets_notouch_[48] ;
 wire \ros_nand4_cap.open_nets_notouch_[49] ;
 wire \ros_nand4_cap.open_nets_notouch_[4] ;
 wire \ros_nand4_cap.open_nets_notouch_[50] ;
 wire \ros_nand4_cap.open_nets_notouch_[51] ;
 wire \ros_nand4_cap.open_nets_notouch_[52] ;
 wire \ros_nand4_cap.open_nets_notouch_[53] ;
 wire \ros_nand4_cap.open_nets_notouch_[54] ;
 wire \ros_nand4_cap.open_nets_notouch_[55] ;
 wire \ros_nand4_cap.open_nets_notouch_[56] ;
 wire \ros_nand4_cap.open_nets_notouch_[57] ;
 wire \ros_nand4_cap.open_nets_notouch_[58] ;
 wire \ros_nand4_cap.open_nets_notouch_[59] ;
 wire \ros_nand4_cap.open_nets_notouch_[5] ;
 wire \ros_nand4_cap.open_nets_notouch_[60] ;
 wire \ros_nand4_cap.open_nets_notouch_[61] ;
 wire \ros_nand4_cap.open_nets_notouch_[62] ;
 wire \ros_nand4_cap.open_nets_notouch_[63] ;
 wire \ros_nand4_cap.open_nets_notouch_[64] ;
 wire \ros_nand4_cap.open_nets_notouch_[65] ;
 wire \ros_nand4_cap.open_nets_notouch_[66] ;
 wire \ros_nand4_cap.open_nets_notouch_[67] ;
 wire \ros_nand4_cap.open_nets_notouch_[68] ;
 wire \ros_nand4_cap.open_nets_notouch_[69] ;
 wire \ros_nand4_cap.open_nets_notouch_[6] ;
 wire \ros_nand4_cap.open_nets_notouch_[70] ;
 wire \ros_nand4_cap.open_nets_notouch_[71] ;
 wire \ros_nand4_cap.open_nets_notouch_[72] ;
 wire \ros_nand4_cap.open_nets_notouch_[73] ;
 wire \ros_nand4_cap.open_nets_notouch_[74] ;
 wire \ros_nand4_cap.open_nets_notouch_[75] ;
 wire \ros_nand4_cap.open_nets_notouch_[76] ;
 wire \ros_nand4_cap.open_nets_notouch_[77] ;
 wire \ros_nand4_cap.open_nets_notouch_[78] ;
 wire \ros_nand4_cap.open_nets_notouch_[79] ;
 wire \ros_nand4_cap.open_nets_notouch_[7] ;
 wire \ros_nand4_cap.open_nets_notouch_[80] ;
 wire \ros_nand4_cap.open_nets_notouch_[81] ;
 wire \ros_nand4_cap.open_nets_notouch_[82] ;
 wire \ros_nand4_cap.open_nets_notouch_[83] ;
 wire \ros_nand4_cap.open_nets_notouch_[84] ;
 wire \ros_nand4_cap.open_nets_notouch_[85] ;
 wire \ros_nand4_cap.open_nets_notouch_[86] ;
 wire \ros_nand4_cap.open_nets_notouch_[87] ;
 wire \ros_nand4_cap.open_nets_notouch_[88] ;
 wire \ros_nand4_cap.open_nets_notouch_[89] ;
 wire \ros_nand4_cap.open_nets_notouch_[8] ;
 wire \ros_nand4_cap.open_nets_notouch_[90] ;
 wire \ros_nand4_cap.open_nets_notouch_[91] ;
 wire \ros_nand4_cap.open_nets_notouch_[92] ;
 wire \ros_nand4_cap.open_nets_notouch_[93] ;
 wire \ros_nand4_cap.open_nets_notouch_[94] ;
 wire \ros_nand4_cap.open_nets_notouch_[95] ;
 wire \ros_nand4_cap.open_nets_notouch_[96] ;
 wire \ros_nand4_cap.open_nets_notouch_[97] ;
 wire \ros_nand4_cap.open_nets_notouch_[98] ;
 wire \ros_nand4_cap.open_nets_notouch_[99] ;
 wire \ros_nand4_cap.open_nets_notouch_[9] ;
 wire \send_counter_syncs[0] ;
 wire \send_counter_syncs[1] ;
 wire \send_counter_syncs[2] ;
 wire \shift_register[0] ;
 wire \shift_register[10] ;
 wire \shift_register[11] ;
 wire \shift_register[12] ;
 wire \shift_register[13] ;
 wire \shift_register[14] ;
 wire \shift_register[15] ;
 wire \shift_register[16] ;
 wire \shift_register[17] ;
 wire \shift_register[18] ;
 wire \shift_register[19] ;
 wire \shift_register[1] ;
 wire \shift_register[20] ;
 wire \shift_register[21] ;
 wire \shift_register[22] ;
 wire \shift_register[23] ;
 wire \shift_register[2] ;
 wire \shift_register[3] ;
 wire \shift_register[4] ;
 wire \shift_register[5] ;
 wire \shift_register[6] ;
 wire \shift_register[7] ;
 wire \shift_register[8] ;
 wire \shift_register[9] ;

 sky130_fd_sc_hd__decap_4 FILLER_0_0_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_257 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_284 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_296 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_95 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_335 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_122 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_154 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_168 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_331 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_138 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_22 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_297 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_295 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_151 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_185 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_74 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_161 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_25 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_318 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_116 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_128 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_140 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_152 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_290 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_302 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_314 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_287 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_313 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_66 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_297 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_144 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_55 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_96 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_291 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_151 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_163 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_175 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_49 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_99 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_332 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_118 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_154 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_329 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_72 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_132 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_44 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_67 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_106 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_318 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_50 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_124 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_70 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_128 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_33 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_36 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_180 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_322 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_334 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_189 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_201 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_324 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_74 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_86 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_100 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_214 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_331 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_35 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_88 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_216 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_129 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__and4_1 _0838_ (.A(\fmeasurment_einv_sub_ros.counts[3] ),
    .B(\fmeasurment_einv_sub_ros.counts[2] ),
    .C(\fmeasurment_einv_sub_ros.counts[1] ),
    .D(\fmeasurment_einv_sub_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _0839_ (.A(\fmeasurment_einv_sub_ros.counts[6] ),
    .B(\fmeasurment_einv_sub_ros.counts[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__and4_1 _0840_ (.A(\fmeasurment_einv_sub_ros.counts[7] ),
    .B(\fmeasurment_einv_sub_ros.counts[4] ),
    .C(_0282_),
    .D(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _0841_ (.A(\fmeasurment_einv_sub_ros.counts[10] ),
    .B(\fmeasurment_einv_sub_ros.counts[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__and4_1 _0842_ (.A(\fmeasurment_einv_sub_ros.counts[11] ),
    .B(\fmeasurment_einv_sub_ros.counts[8] ),
    .C(_0284_),
    .D(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_2 _0843_ (.A(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__and4_1 _0844_ (.A(\fmeasurment_einv_sub_ros.counts[14] ),
    .B(\fmeasurment_einv_sub_ros.counts[13] ),
    .C(\fmeasurment_einv_sub_ros.counts[12] ),
    .D(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_2 _0845_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__and4_2 _0846_ (.A(\fmeasurment_einv_sub_ros.counts[17] ),
    .B(\fmeasurment_einv_sub_ros.counts[16] ),
    .C(\fmeasurment_einv_sub_ros.counts[15] ),
    .D(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__a21oi_1 _0847_ (.A1(\fmeasurment_einv_sub_ros.counts[18] ),
    .A2(_0290_),
    .B1(\fmeasurment_einv_sub_ros.counts[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0291_));
 sky130_fd_sc_hd__buf_2 _0848_ (.A(\fmeasurment_einv_sub_ros.reset_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__a31o_1 _0849_ (.A1(\fmeasurment_einv_sub_ros.counts[19] ),
    .A2(\fmeasurment_einv_sub_ros.counts[18] ),
    .A3(_0290_),
    .B1(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(_0291_),
    .B(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0281_));
 sky130_fd_sc_hd__clkbuf_4 _0851_ (.A(\fmeasurment_einv_sub_ros.reset_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__a21oi_1 _0852_ (.A1(\fmeasurment_einv_sub_ros.counts[18] ),
    .A2(_0290_),
    .B1(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0295_));
 sky130_fd_sc_hd__o21a_1 _0853_ (.A1(\fmeasurment_einv_sub_ros.counts[18] ),
    .A2(_0290_),
    .B1(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__and3_1 _0854_ (.A(\fmeasurment_einv_sub_ros.counts[16] ),
    .B(\fmeasurment_einv_sub_ros.counts[15] ),
    .C(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(_0294_),
    .B(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0297_));
 sky130_fd_sc_hd__o21a_1 _0856_ (.A1(\fmeasurment_einv_sub_ros.counts[17] ),
    .A2(_0296_),
    .B1(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _0857_ (.A1(\fmeasurment_einv_sub_ros.counts[15] ),
    .A2(_0289_),
    .B1(\fmeasurment_einv_sub_ros.counts[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0298_));
 sky130_fd_sc_hd__nor3_1 _0858_ (.A(_0294_),
    .B(_0296_),
    .C(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0278_));
 sky130_fd_sc_hd__a21oi_1 _0859_ (.A1(\fmeasurment_einv_sub_ros.counts[15] ),
    .A2(_0289_),
    .B1(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0299_));
 sky130_fd_sc_hd__o21a_1 _0860_ (.A1(\fmeasurment_einv_sub_ros.counts[15] ),
    .A2(_0289_),
    .B1(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__and3_1 _0861_ (.A(\fmeasurment_einv_sub_ros.counts[13] ),
    .B(\fmeasurment_einv_sub_ros.counts[12] ),
    .C(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__nor2_1 _0862_ (.A(_0294_),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0301_));
 sky130_fd_sc_hd__o21a_1 _0863_ (.A1(\fmeasurment_einv_sub_ros.counts[14] ),
    .A2(_0300_),
    .B1(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__a21oi_1 _0864_ (.A1(\fmeasurment_einv_sub_ros.counts[12] ),
    .A2(_0287_),
    .B1(\fmeasurment_einv_sub_ros.counts[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0302_));
 sky130_fd_sc_hd__nor3_1 _0865_ (.A(_0294_),
    .B(_0300_),
    .C(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0275_));
 sky130_fd_sc_hd__a21oi_1 _0866_ (.A1(\fmeasurment_einv_sub_ros.counts[12] ),
    .A2(_0287_),
    .B1(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0303_));
 sky130_fd_sc_hd__o21a_1 _0867_ (.A1(\fmeasurment_einv_sub_ros.counts[12] ),
    .A2(_0287_),
    .B1(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__and3_1 _0868_ (.A(\fmeasurment_einv_sub_ros.counts[8] ),
    .B(_0284_),
    .C(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__nor2_1 _0869_ (.A(_0292_),
    .B(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0305_));
 sky130_fd_sc_hd__o21a_1 _0870_ (.A1(\fmeasurment_einv_sub_ros.counts[11] ),
    .A2(_0304_),
    .B1(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__and3_1 _0871_ (.A(\fmeasurment_einv_sub_ros.counts[9] ),
    .B(\fmeasurment_einv_sub_ros.counts[8] ),
    .C(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__nor2_1 _0872_ (.A(_0292_),
    .B(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0307_));
 sky130_fd_sc_hd__o21a_1 _0873_ (.A1(\fmeasurment_einv_sub_ros.counts[10] ),
    .A2(_0306_),
    .B1(_0307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _0874_ (.A(\fmeasurment_einv_sub_ros.counts[8] ),
    .B(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _0875_ (.A(_0292_),
    .B(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0309_));
 sky130_fd_sc_hd__o21a_1 _0876_ (.A1(\fmeasurment_einv_sub_ros.counts[9] ),
    .A2(_0308_),
    .B1(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(_0292_),
    .B(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0310_));
 sky130_fd_sc_hd__o21a_1 _0878_ (.A1(\fmeasurment_einv_sub_ros.counts[8] ),
    .A2(_0284_),
    .B1(_0310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _0879_ (.A(\fmeasurment_einv_sub_ros.counts[4] ),
    .B(_0282_),
    .C(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _0880_ (.A(_0292_),
    .B(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0312_));
 sky130_fd_sc_hd__o21a_1 _0881_ (.A1(\fmeasurment_einv_sub_ros.counts[7] ),
    .A2(_0311_),
    .B1(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__and3_1 _0882_ (.A(\fmeasurment_einv_sub_ros.counts[5] ),
    .B(\fmeasurment_einv_sub_ros.counts[4] ),
    .C(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__nor2_1 _0883_ (.A(_0292_),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0314_));
 sky130_fd_sc_hd__o21a_1 _0884_ (.A1(\fmeasurment_einv_sub_ros.counts[6] ),
    .A2(_0313_),
    .B1(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0268_));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(\fmeasurment_einv_sub_ros.counts[4] ),
    .B(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__nor2_1 _0886_ (.A(_0292_),
    .B(_0313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0316_));
 sky130_fd_sc_hd__o21a_1 _0887_ (.A1(\fmeasurment_einv_sub_ros.counts[5] ),
    .A2(_0315_),
    .B1(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_1 _0888_ (.A(_0292_),
    .B(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0317_));
 sky130_fd_sc_hd__o21a_1 _0889_ (.A1(\fmeasurment_einv_sub_ros.counts[4] ),
    .A2(_0282_),
    .B1(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _0890_ (.A(\fmeasurment_einv_sub_ros.counts[2] ),
    .B(\fmeasurment_einv_sub_ros.counts[1] ),
    .C(\fmeasurment_einv_sub_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_1 _0891_ (.A(_0292_),
    .B(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0319_));
 sky130_fd_sc_hd__o21a_1 _0892_ (.A1(\fmeasurment_einv_sub_ros.counts[3] ),
    .A2(_0318_),
    .B1(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _0893_ (.A1(\fmeasurment_einv_sub_ros.counts[1] ),
    .A2(\fmeasurment_einv_sub_ros.counts[0] ),
    .B1(\fmeasurment_einv_sub_ros.counts[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0320_));
 sky130_fd_sc_hd__nor3_1 _0894_ (.A(_0294_),
    .B(_0318_),
    .C(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0264_));
 sky130_fd_sc_hd__a21oi_1 _0895_ (.A1(\fmeasurment_einv_sub_ros.counts[1] ),
    .A2(\fmeasurment_einv_sub_ros.counts[0] ),
    .B1(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0321_));
 sky130_fd_sc_hd__o21a_1 _0896_ (.A1(\fmeasurment_einv_sub_ros.counts[1] ),
    .A2(\fmeasurment_einv_sub_ros.counts[0] ),
    .B1(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(_0294_),
    .B(\fmeasurment_einv_sub_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0262_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(net2),
    .A1(\fmeasurment_einv_sub_ros.latch_counter_syncs[2] ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_4 _0899_ (.A(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[19] ),
    .A1(\fmeasurment_einv_sub_ros.counts[19] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[18] ),
    .A1(\fmeasurment_einv_sub_ros.counts[18] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _0903_ (.A(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[17] ),
    .A1(\fmeasurment_einv_sub_ros.counts[17] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0905_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[16] ),
    .A1(\fmeasurment_einv_sub_ros.counts[16] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0907_ (.A(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[15] ),
    .A1(\fmeasurment_einv_sub_ros.counts[15] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0909_ (.A(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[14] ),
    .A1(\fmeasurment_einv_sub_ros.counts[14] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[13] ),
    .A1(\fmeasurment_einv_sub_ros.counts[13] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0913_ (.A(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[12] ),
    .A1(\fmeasurment_einv_sub_ros.counts[12] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _0915_ (.A(_0331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[11] ),
    .A1(\fmeasurment_einv_sub_ros.counts[11] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0917_ (.A(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[10] ),
    .A1(\fmeasurment_einv_sub_ros.counts[10] ),
    .S(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _0919_ (.A(_0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__buf_4 _0920_ (.A(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _0921_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[9] ),
    .A1(\fmeasurment_einv_sub_ros.counts[9] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0922_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0923_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[8] ),
    .A1(\fmeasurment_einv_sub_ros.counts[8] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _0924_ (.A(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _0925_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[7] ),
    .A1(\fmeasurment_einv_sub_ros.counts[7] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _0926_ (.A(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[6] ),
    .A1(\fmeasurment_einv_sub_ros.counts[6] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _0928_ (.A(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[5] ),
    .A1(\fmeasurment_einv_sub_ros.counts[5] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0930_ (.A(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[4] ),
    .A1(\fmeasurment_einv_sub_ros.counts[4] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0932_ (.A(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[3] ),
    .A1(\fmeasurment_einv_sub_ros.counts[3] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0934_ (.A(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[2] ),
    .A1(\fmeasurment_einv_sub_ros.counts[2] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _0936_ (.A(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[1] ),
    .A1(\fmeasurment_einv_sub_ros.counts[1] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _0938_ (.A(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(\fmeasurment_einv_sub_ros.cycle_count[0] ),
    .A1(\fmeasurment_einv_sub_ros.counts[0] ),
    .S(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0940_ (.A(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__and4_1 _0941_ (.A(\fmeasurment_nand4_cap_ros.counts[3] ),
    .B(\fmeasurment_nand4_cap_ros.counts[2] ),
    .C(\fmeasurment_nand4_cap_ros.counts[1] ),
    .D(\fmeasurment_nand4_cap_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__and2_1 _0942_ (.A(\fmeasurment_nand4_cap_ros.counts[6] ),
    .B(\fmeasurment_nand4_cap_ros.counts[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__and4_1 _0943_ (.A(\fmeasurment_nand4_cap_ros.counts[7] ),
    .B(\fmeasurment_nand4_cap_ros.counts[4] ),
    .C(_0345_),
    .D(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__and2_1 _0944_ (.A(\fmeasurment_nand4_cap_ros.counts[10] ),
    .B(\fmeasurment_nand4_cap_ros.counts[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__and4_1 _0945_ (.A(\fmeasurment_nand4_cap_ros.counts[11] ),
    .B(\fmeasurment_nand4_cap_ros.counts[8] ),
    .C(_0347_),
    .D(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0946_ (.A(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__and4_1 _0947_ (.A(\fmeasurment_nand4_cap_ros.counts[14] ),
    .B(\fmeasurment_nand4_cap_ros.counts[13] ),
    .C(\fmeasurment_nand4_cap_ros.counts[12] ),
    .D(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_2 _0948_ (.A(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__and4_1 _0949_ (.A(\fmeasurment_nand4_cap_ros.counts[17] ),
    .B(\fmeasurment_nand4_cap_ros.counts[16] ),
    .C(\fmeasurment_nand4_cap_ros.counts[15] ),
    .D(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__a21oi_1 _0950_ (.A1(\fmeasurment_nand4_cap_ros.counts[18] ),
    .A2(_0353_),
    .B1(\fmeasurment_nand4_cap_ros.counts[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0354_));
 sky130_fd_sc_hd__buf_2 _0951_ (.A(\fmeasurment_nand4_cap_ros.reset_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__a31o_1 _0952_ (.A1(\fmeasurment_nand4_cap_ros.counts[19] ),
    .A2(\fmeasurment_nand4_cap_ros.counts[18] ),
    .A3(_0353_),
    .B1(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__nor2_1 _0953_ (.A(_0354_),
    .B(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0241_));
 sky130_fd_sc_hd__clkbuf_4 _0954_ (.A(\fmeasurment_nand4_cap_ros.reset_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__a21oi_1 _0955_ (.A1(\fmeasurment_nand4_cap_ros.counts[18] ),
    .A2(_0353_),
    .B1(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0358_));
 sky130_fd_sc_hd__o21a_1 _0956_ (.A1(\fmeasurment_nand4_cap_ros.counts[18] ),
    .A2(_0353_),
    .B1(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__and3_1 _0957_ (.A(\fmeasurment_nand4_cap_ros.counts[16] ),
    .B(\fmeasurment_nand4_cap_ros.counts[15] ),
    .C(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _0958_ (.A(_0357_),
    .B(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0360_));
 sky130_fd_sc_hd__o21a_1 _0959_ (.A1(\fmeasurment_nand4_cap_ros.counts[17] ),
    .A2(_0359_),
    .B1(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__a21oi_1 _0960_ (.A1(\fmeasurment_nand4_cap_ros.counts[15] ),
    .A2(_0352_),
    .B1(\fmeasurment_nand4_cap_ros.counts[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0361_));
 sky130_fd_sc_hd__nor3_1 _0961_ (.A(_0357_),
    .B(_0359_),
    .C(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0238_));
 sky130_fd_sc_hd__a21oi_1 _0962_ (.A1(\fmeasurment_nand4_cap_ros.counts[15] ),
    .A2(_0352_),
    .B1(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0362_));
 sky130_fd_sc_hd__o21a_1 _0963_ (.A1(\fmeasurment_nand4_cap_ros.counts[15] ),
    .A2(_0352_),
    .B1(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__and3_1 _0964_ (.A(\fmeasurment_nand4_cap_ros.counts[13] ),
    .B(\fmeasurment_nand4_cap_ros.counts[12] ),
    .C(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_1 _0965_ (.A(_0357_),
    .B(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0364_));
 sky130_fd_sc_hd__o21a_1 _0966_ (.A1(\fmeasurment_nand4_cap_ros.counts[14] ),
    .A2(_0363_),
    .B1(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__a21oi_1 _0967_ (.A1(\fmeasurment_nand4_cap_ros.counts[12] ),
    .A2(_0350_),
    .B1(\fmeasurment_nand4_cap_ros.counts[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0365_));
 sky130_fd_sc_hd__nor3_1 _0968_ (.A(_0357_),
    .B(_0363_),
    .C(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0235_));
 sky130_fd_sc_hd__a21oi_1 _0969_ (.A1(\fmeasurment_nand4_cap_ros.counts[12] ),
    .A2(_0350_),
    .B1(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0366_));
 sky130_fd_sc_hd__o21a_1 _0970_ (.A1(\fmeasurment_nand4_cap_ros.counts[12] ),
    .A2(_0350_),
    .B1(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0234_));
 sky130_fd_sc_hd__and3_1 _0971_ (.A(\fmeasurment_nand4_cap_ros.counts[8] ),
    .B(_0347_),
    .C(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__nor2_1 _0972_ (.A(_0355_),
    .B(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0368_));
 sky130_fd_sc_hd__o21a_1 _0973_ (.A1(\fmeasurment_nand4_cap_ros.counts[11] ),
    .A2(_0367_),
    .B1(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__and3_1 _0974_ (.A(\fmeasurment_nand4_cap_ros.counts[9] ),
    .B(\fmeasurment_nand4_cap_ros.counts[8] ),
    .C(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__nor2_1 _0975_ (.A(_0355_),
    .B(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0370_));
 sky130_fd_sc_hd__o21a_1 _0976_ (.A1(\fmeasurment_nand4_cap_ros.counts[10] ),
    .A2(_0369_),
    .B1(_0370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__and2_1 _0977_ (.A(\fmeasurment_nand4_cap_ros.counts[8] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _0978_ (.A(_0355_),
    .B(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0372_));
 sky130_fd_sc_hd__o21a_1 _0979_ (.A1(\fmeasurment_nand4_cap_ros.counts[9] ),
    .A2(_0371_),
    .B1(_0372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _0980_ (.A(_0355_),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0373_));
 sky130_fd_sc_hd__o21a_1 _0981_ (.A1(\fmeasurment_nand4_cap_ros.counts[8] ),
    .A2(_0347_),
    .B1(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__and3_1 _0982_ (.A(\fmeasurment_nand4_cap_ros.counts[4] ),
    .B(_0345_),
    .C(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_1 _0983_ (.A(_0355_),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0375_));
 sky130_fd_sc_hd__o21a_1 _0984_ (.A1(\fmeasurment_nand4_cap_ros.counts[7] ),
    .A2(_0374_),
    .B1(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0229_));
 sky130_fd_sc_hd__and3_1 _0985_ (.A(\fmeasurment_nand4_cap_ros.counts[5] ),
    .B(\fmeasurment_nand4_cap_ros.counts[4] ),
    .C(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_1 _0986_ (.A(_0355_),
    .B(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0377_));
 sky130_fd_sc_hd__o21a_1 _0987_ (.A1(\fmeasurment_nand4_cap_ros.counts[6] ),
    .A2(_0376_),
    .B1(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _0988_ (.A(\fmeasurment_nand4_cap_ros.counts[4] ),
    .B(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(_0355_),
    .B(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0379_));
 sky130_fd_sc_hd__o21a_1 _0990_ (.A1(\fmeasurment_nand4_cap_ros.counts[5] ),
    .A2(_0378_),
    .B1(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _0991_ (.A(_0355_),
    .B(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0380_));
 sky130_fd_sc_hd__o21a_1 _0992_ (.A1(\fmeasurment_nand4_cap_ros.counts[4] ),
    .A2(_0345_),
    .B1(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0226_));
 sky130_fd_sc_hd__and3_1 _0993_ (.A(\fmeasurment_nand4_cap_ros.counts[2] ),
    .B(\fmeasurment_nand4_cap_ros.counts[1] ),
    .C(\fmeasurment_nand4_cap_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__nor2_1 _0994_ (.A(_0355_),
    .B(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0382_));
 sky130_fd_sc_hd__o21a_1 _0995_ (.A1(\fmeasurment_nand4_cap_ros.counts[3] ),
    .A2(_0381_),
    .B1(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__a21oi_1 _0996_ (.A1(\fmeasurment_nand4_cap_ros.counts[1] ),
    .A2(\fmeasurment_nand4_cap_ros.counts[0] ),
    .B1(\fmeasurment_nand4_cap_ros.counts[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0383_));
 sky130_fd_sc_hd__nor3_1 _0997_ (.A(_0357_),
    .B(_0381_),
    .C(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0224_));
 sky130_fd_sc_hd__a21oi_1 _0998_ (.A1(\fmeasurment_nand4_cap_ros.counts[1] ),
    .A2(\fmeasurment_nand4_cap_ros.counts[0] ),
    .B1(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0384_));
 sky130_fd_sc_hd__o21a_1 _0999_ (.A1(\fmeasurment_nand4_cap_ros.counts[1] ),
    .A2(\fmeasurment_nand4_cap_ros.counts[0] ),
    .B1(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _1000_ (.A(_0357_),
    .B(\fmeasurment_nand4_cap_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0222_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(net2),
    .A1(\fmeasurment_nand4_ros.latch_counter_syncs[2] ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_4 _1002_ (.A(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(\fmeasurment_nand4_ros.cycle_count[19] ),
    .A1(\fmeasurment_nand4_ros.counts[19] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(\fmeasurment_nand4_ros.cycle_count[18] ),
    .A1(\fmeasurment_nand4_ros.counts[18] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(\fmeasurment_nand4_ros.cycle_count[17] ),
    .A1(\fmeasurment_nand4_ros.counts[17] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _1008_ (.A(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1009_ (.A0(\fmeasurment_nand4_ros.cycle_count[16] ),
    .A1(\fmeasurment_nand4_ros.counts[16] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _1010_ (.A(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(\fmeasurment_nand4_ros.cycle_count[15] ),
    .A1(\fmeasurment_nand4_ros.counts[15] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(\fmeasurment_nand4_ros.cycle_count[14] ),
    .A1(\fmeasurment_nand4_ros.counts[14] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _1014_ (.A(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1015_ (.A0(\fmeasurment_nand4_ros.cycle_count[13] ),
    .A1(\fmeasurment_nand4_ros.counts[13] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _1016_ (.A(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1017_ (.A0(\fmeasurment_nand4_ros.cycle_count[12] ),
    .A1(\fmeasurment_nand4_ros.counts[12] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _1018_ (.A(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(\fmeasurment_nand4_ros.cycle_count[11] ),
    .A1(\fmeasurment_nand4_ros.counts[11] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _1020_ (.A(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(\fmeasurment_nand4_ros.cycle_count[10] ),
    .A1(\fmeasurment_nand4_ros.counts[10] ),
    .S(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_4 _1023_ (.A(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(\fmeasurment_nand4_ros.cycle_count[9] ),
    .A1(\fmeasurment_nand4_ros.counts[9] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1026_ (.A0(\fmeasurment_nand4_ros.cycle_count[8] ),
    .A1(\fmeasurment_nand4_ros.counts[8] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _1027_ (.A(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(\fmeasurment_nand4_ros.cycle_count[7] ),
    .A1(\fmeasurment_nand4_ros.counts[7] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _1029_ (.A(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\fmeasurment_nand4_ros.cycle_count[6] ),
    .A1(\fmeasurment_nand4_ros.counts[6] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(\fmeasurment_nand4_ros.cycle_count[5] ),
    .A1(\fmeasurment_nand4_ros.counts[5] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _1033_ (.A(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(\fmeasurment_nand4_ros.cycle_count[4] ),
    .A1(\fmeasurment_nand4_ros.counts[4] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _1035_ (.A(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _1036_ (.A0(\fmeasurment_nand4_ros.cycle_count[3] ),
    .A1(\fmeasurment_nand4_ros.counts[3] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _1037_ (.A(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1038_ (.A0(\fmeasurment_nand4_ros.cycle_count[2] ),
    .A1(\fmeasurment_nand4_ros.counts[2] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _1039_ (.A(_0405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(\fmeasurment_nand4_ros.cycle_count[1] ),
    .A1(\fmeasurment_nand4_ros.counts[1] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _1042_ (.A0(\fmeasurment_nand4_ros.cycle_count[0] ),
    .A1(\fmeasurment_nand4_ros.counts[0] ),
    .S(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _1043_ (.A(_0407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(net2),
    .A1(\fmeasurment_nand4_cap_ros.latch_counter_syncs[2] ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_4 _1045_ (.A(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[19] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[19] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _1048_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[18] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[18] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _1049_ (.A(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[17] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[17] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[16] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[16] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[15] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[15] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[14] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[14] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _1057_ (.A(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1058_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[13] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[13] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _1059_ (.A(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _1060_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[12] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[12] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _1062_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[11] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[11] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1063_ (.A(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[10] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[10] ),
    .S(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1065_ (.A(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _1066_ (.A(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _1067_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[9] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[9] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1068_ (.A(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _1069_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[8] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[8] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1070_ (.A(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _1071_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[7] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[7] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _1072_ (.A(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _1073_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[6] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[6] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _1075_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[5] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[5] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _1076_ (.A(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _1077_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[4] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[4] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _1079_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[3] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[3] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _1080_ (.A(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _1081_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[2] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[2] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _1082_ (.A(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _1083_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[1] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[1] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _1084_ (.A(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _1085_ (.A0(\fmeasurment_nand4_cap_ros.cycle_count[0] ),
    .A1(\fmeasurment_nand4_cap_ros.counts[0] ),
    .S(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1086_ (.A(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__and4_1 _1087_ (.A(\fmeasurment_nand4_ros.counts[3] ),
    .B(\fmeasurment_nand4_ros.counts[2] ),
    .C(\fmeasurment_nand4_ros.counts[1] ),
    .D(\fmeasurment_nand4_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _1088_ (.A(\fmeasurment_nand4_ros.counts[6] ),
    .B(\fmeasurment_nand4_ros.counts[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__and4_1 _1089_ (.A(\fmeasurment_nand4_ros.counts[7] ),
    .B(\fmeasurment_nand4_ros.counts[4] ),
    .C(_0431_),
    .D(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _1090_ (.A(\fmeasurment_nand4_ros.counts[10] ),
    .B(\fmeasurment_nand4_ros.counts[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__and4_1 _1091_ (.A(\fmeasurment_nand4_ros.counts[11] ),
    .B(\fmeasurment_nand4_ros.counts[8] ),
    .C(_0433_),
    .D(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1092_ (.A(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__and4_1 _1093_ (.A(\fmeasurment_nand4_ros.counts[14] ),
    .B(\fmeasurment_nand4_ros.counts[13] ),
    .C(\fmeasurment_nand4_ros.counts[12] ),
    .D(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0437_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1094_ (.A(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__and4_1 _1095_ (.A(\fmeasurment_nand4_ros.counts[17] ),
    .B(\fmeasurment_nand4_ros.counts[16] ),
    .C(\fmeasurment_nand4_ros.counts[15] ),
    .D(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1096_ (.A1(\fmeasurment_nand4_ros.counts[18] ),
    .A2(_0439_),
    .B1(\fmeasurment_nand4_ros.counts[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0440_));
 sky130_fd_sc_hd__buf_2 _1097_ (.A(\fmeasurment_nand4_ros.reset_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0441_));
 sky130_fd_sc_hd__a31o_1 _1098_ (.A1(\fmeasurment_nand4_ros.counts[19] ),
    .A2(\fmeasurment_nand4_ros.counts[18] ),
    .A3(_0439_),
    .B1(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_1 _1099_ (.A(_0440_),
    .B(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0181_));
 sky130_fd_sc_hd__clkbuf_4 _1100_ (.A(\fmeasurment_nand4_ros.reset_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__a21oi_1 _1101_ (.A1(\fmeasurment_nand4_ros.counts[18] ),
    .A2(_0439_),
    .B1(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0444_));
 sky130_fd_sc_hd__o21a_1 _1102_ (.A1(\fmeasurment_nand4_ros.counts[18] ),
    .A2(_0439_),
    .B1(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__and3_1 _1103_ (.A(\fmeasurment_nand4_ros.counts[16] ),
    .B(\fmeasurment_nand4_ros.counts[15] ),
    .C(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_1 _1104_ (.A(_0443_),
    .B(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0446_));
 sky130_fd_sc_hd__o21a_1 _1105_ (.A1(\fmeasurment_nand4_ros.counts[17] ),
    .A2(_0445_),
    .B1(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__a21oi_1 _1106_ (.A1(\fmeasurment_nand4_ros.counts[15] ),
    .A2(_0438_),
    .B1(\fmeasurment_nand4_ros.counts[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0447_));
 sky130_fd_sc_hd__nor3_1 _1107_ (.A(_0443_),
    .B(_0445_),
    .C(_0447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0178_));
 sky130_fd_sc_hd__a21oi_1 _1108_ (.A1(\fmeasurment_nand4_ros.counts[15] ),
    .A2(_0438_),
    .B1(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0448_));
 sky130_fd_sc_hd__o21a_1 _1109_ (.A1(\fmeasurment_nand4_ros.counts[15] ),
    .A2(_0438_),
    .B1(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _1110_ (.A(\fmeasurment_nand4_ros.counts[13] ),
    .B(\fmeasurment_nand4_ros.counts[12] ),
    .C(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__nor2_1 _1111_ (.A(_0443_),
    .B(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0450_));
 sky130_fd_sc_hd__o21a_1 _1112_ (.A1(\fmeasurment_nand4_ros.counts[14] ),
    .A2(_0449_),
    .B1(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__a21oi_1 _1113_ (.A1(\fmeasurment_nand4_ros.counts[12] ),
    .A2(_0436_),
    .B1(\fmeasurment_nand4_ros.counts[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0451_));
 sky130_fd_sc_hd__nor3_1 _1114_ (.A(_0443_),
    .B(_0449_),
    .C(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0175_));
 sky130_fd_sc_hd__a21oi_1 _1115_ (.A1(\fmeasurment_nand4_ros.counts[12] ),
    .A2(_0436_),
    .B1(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0452_));
 sky130_fd_sc_hd__o21a_1 _1116_ (.A1(\fmeasurment_nand4_ros.counts[12] ),
    .A2(_0436_),
    .B1(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__and3_1 _1117_ (.A(\fmeasurment_nand4_ros.counts[8] ),
    .B(_0433_),
    .C(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _1118_ (.A(_0441_),
    .B(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0454_));
 sky130_fd_sc_hd__o21a_1 _1119_ (.A1(\fmeasurment_nand4_ros.counts[11] ),
    .A2(_0453_),
    .B1(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__and3_1 _1120_ (.A(\fmeasurment_nand4_ros.counts[9] ),
    .B(\fmeasurment_nand4_ros.counts[8] ),
    .C(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _1121_ (.A(_0441_),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0456_));
 sky130_fd_sc_hd__o21a_1 _1122_ (.A1(\fmeasurment_nand4_ros.counts[10] ),
    .A2(_0455_),
    .B1(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _1123_ (.A(\fmeasurment_nand4_ros.counts[8] ),
    .B(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0457_));
 sky130_fd_sc_hd__nor2_1 _1124_ (.A(_0441_),
    .B(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0458_));
 sky130_fd_sc_hd__o21a_1 _1125_ (.A1(\fmeasurment_nand4_ros.counts[9] ),
    .A2(_0457_),
    .B1(_0458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _1126_ (.A(_0441_),
    .B(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0459_));
 sky130_fd_sc_hd__o21a_1 _1127_ (.A1(\fmeasurment_nand4_ros.counts[8] ),
    .A2(_0433_),
    .B1(_0459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__and3_1 _1128_ (.A(\fmeasurment_nand4_ros.counts[4] ),
    .B(_0431_),
    .C(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _1129_ (.A(_0441_),
    .B(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0461_));
 sky130_fd_sc_hd__o21a_1 _1130_ (.A1(\fmeasurment_nand4_ros.counts[7] ),
    .A2(_0460_),
    .B1(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__and3_1 _1131_ (.A(\fmeasurment_nand4_ros.counts[5] ),
    .B(\fmeasurment_nand4_ros.counts[4] ),
    .C(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0462_));
 sky130_fd_sc_hd__nor2_1 _1132_ (.A(_0441_),
    .B(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0463_));
 sky130_fd_sc_hd__o21a_1 _1133_ (.A1(\fmeasurment_nand4_ros.counts[6] ),
    .A2(_0462_),
    .B1(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _1134_ (.A(\fmeasurment_nand4_ros.counts[4] ),
    .B(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _1135_ (.A(_0441_),
    .B(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_1 _1136_ (.A1(\fmeasurment_nand4_ros.counts[5] ),
    .A2(_0464_),
    .B1(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__nor2_1 _1137_ (.A(_0441_),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0466_));
 sky130_fd_sc_hd__o21a_1 _1138_ (.A1(\fmeasurment_nand4_ros.counts[4] ),
    .A2(_0431_),
    .B1(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__and3_1 _1139_ (.A(\fmeasurment_nand4_ros.counts[2] ),
    .B(\fmeasurment_nand4_ros.counts[1] ),
    .C(\fmeasurment_nand4_ros.counts[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0467_));
 sky130_fd_sc_hd__nor2_1 _1140_ (.A(_0441_),
    .B(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0468_));
 sky130_fd_sc_hd__o21a_1 _1141_ (.A1(\fmeasurment_nand4_ros.counts[3] ),
    .A2(_0467_),
    .B1(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__a21oi_1 _1142_ (.A1(\fmeasurment_nand4_ros.counts[1] ),
    .A2(\fmeasurment_nand4_ros.counts[0] ),
    .B1(\fmeasurment_nand4_ros.counts[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0469_));
 sky130_fd_sc_hd__nor3_1 _1143_ (.A(_0443_),
    .B(_0467_),
    .C(_0469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0164_));
 sky130_fd_sc_hd__a21oi_1 _1144_ (.A1(\fmeasurment_nand4_ros.counts[1] ),
    .A2(\fmeasurment_nand4_ros.counts[0] ),
    .B1(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0470_));
 sky130_fd_sc_hd__o21a_1 _1145_ (.A1(\fmeasurment_nand4_ros.counts[1] ),
    .A2(\fmeasurment_nand4_ros.counts[0] ),
    .B1(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_1 _1146_ (.A(\fmeasurment_nand4_ros.counts[0] ),
    .B(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0162_));
 sky130_fd_sc_hd__or2_1 _1147_ (.A(net8),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _1148_ (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0472_));
 sky130_fd_sc_hd__nor2_1 _1149_ (.A(_0472_),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0473_));
 sky130_fd_sc_hd__and2_1 _1150_ (.A(\fmeasurment_nand4_ros.counts[3] ),
    .B(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0474_));
 sky130_fd_sc_hd__and3_1 _1151_ (.A(\fmeasurment_nand4_ros.counts[7] ),
    .B(net8),
    .C(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_1 _1152_ (.A(net8),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0476_));
 sky130_fd_sc_hd__a2111o_1 _1153_ (.A1(\fmeasurment_nand4_ros.counts[5] ),
    .A2(_0472_),
    .B1(_0474_),
    .C1(_0475_),
    .D1(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0477_));
 sky130_fd_sc_hd__o21ai_1 _1154_ (.A1(\fmeasurment_nand4_ros.counts[1] ),
    .A2(_0471_),
    .B1(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fmeasurment_nand4_ros.divided_clk ));
 sky130_fd_sc_hd__a221o_1 _1155_ (.A1(\fmeasurment_nand4_cap_ros.counts[5] ),
    .A2(_0472_),
    .B1(_0473_),
    .B2(\fmeasurment_nand4_cap_ros.counts[3] ),
    .C1(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0478_));
 sky130_fd_sc_hd__a31o_1 _1156_ (.A1(\fmeasurment_nand4_cap_ros.counts[7] ),
    .A2(net8),
    .A3(net9),
    .B1(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0479_));
 sky130_fd_sc_hd__o21ai_1 _1157_ (.A1(\fmeasurment_nand4_cap_ros.counts[1] ),
    .A2(_0471_),
    .B1(_0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fmeasurment_nand4_cap_ros.divided_clk ));
 sky130_fd_sc_hd__a221o_1 _1158_ (.A1(\fmeasurment_einv_sub_ros.counts[5] ),
    .A2(_0472_),
    .B1(_0473_),
    .B2(\fmeasurment_einv_sub_ros.counts[3] ),
    .C1(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0480_));
 sky130_fd_sc_hd__a31o_1 _1159_ (.A1(\fmeasurment_einv_sub_ros.counts[7] ),
    .A2(net8),
    .A3(net9),
    .B1(_0480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0481_));
 sky130_fd_sc_hd__o21ai_1 _1160_ (.A1(\fmeasurment_einv_sub_ros.counts[1] ),
    .A2(_0471_),
    .B1(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fmeasurment_einv_sub_ros.divided_clk ));
 sky130_fd_sc_hd__xor2_2 _1161_ (.A(clknet_2_2__leaf_clk),
    .B(\shift_register[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(data_stream));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0482_));
 sky130_fd_sc_hd__buf_2 _1163_ (.A(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0483_));
 sky130_fd_sc_hd__nor2_2 _1164_ (.A(\send_counter_syncs[2] ),
    .B(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0484_));
 sky130_fd_sc_hd__clkbuf_4 _1165_ (.A(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0485_));
 sky130_fd_sc_hd__or2_1 _1166_ (.A(net6),
    .B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0486_));
 sky130_fd_sc_hd__buf_2 _1167_ (.A(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0487_));
 sky130_fd_sc_hd__inv_2 _1168_ (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0489_));
 sky130_fd_sc_hd__o21a_1 _1170_ (.A1(_0488_),
    .A2(_0489_),
    .B1(\send_counter_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0490_));
 sky130_fd_sc_hd__buf_2 _1171_ (.A(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _1172_ (.A(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0492_));
 sky130_fd_sc_hd__buf_2 _1173_ (.A(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0493_));
 sky130_fd_sc_hd__buf_2 _1174_ (.A(\ena_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0494_));
 sky130_fd_sc_hd__o221a_1 _1175_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[1] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[1] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0495_));
 sky130_fd_sc_hd__o211a_1 _1176_ (.A1(\fmeasurment_nand4_ros.cycle_count[1] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0496_));
 sky130_fd_sc_hd__a221o_1 _1177_ (.A1(net318),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net316),
    .C1(_0496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__o221a_1 _1178_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[2] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[2] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0497_));
 sky130_fd_sc_hd__o211a_1 _1179_ (.A1(\fmeasurment_nand4_ros.cycle_count[2] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0498_));
 sky130_fd_sc_hd__a221o_1 _1180_ (.A1(net333),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net318),
    .C1(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__o221a_1 _1181_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[3] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[3] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0499_));
 sky130_fd_sc_hd__o211a_1 _1182_ (.A1(\fmeasurment_nand4_ros.cycle_count[3] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0500_));
 sky130_fd_sc_hd__a221o_1 _1183_ (.A1(net346),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net333),
    .C1(_0500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__o221a_1 _1184_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[4] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[4] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0501_));
 sky130_fd_sc_hd__o211a_1 _1185_ (.A1(\fmeasurment_nand4_ros.cycle_count[4] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0502_));
 sky130_fd_sc_hd__a221o_1 _1186_ (.A1(net340),
    .A2(_0483_),
    .B1(_0485_),
    .B2(\shift_register[3] ),
    .C1(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__o221a_1 _1187_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[5] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[5] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0503_));
 sky130_fd_sc_hd__o211a_1 _1188_ (.A1(\fmeasurment_nand4_ros.cycle_count[5] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0504_));
 sky130_fd_sc_hd__a221o_1 _1189_ (.A1(net330),
    .A2(_0483_),
    .B1(_0485_),
    .B2(\shift_register[4] ),
    .C1(_0504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__o221a_1 _1190_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[6] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[6] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0505_));
 sky130_fd_sc_hd__o211a_1 _1191_ (.A1(\fmeasurment_nand4_ros.cycle_count[6] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0506_));
 sky130_fd_sc_hd__a221o_1 _1192_ (.A1(net334),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net330),
    .C1(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__o221a_1 _1193_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[7] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[7] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0507_));
 sky130_fd_sc_hd__o211a_1 _1194_ (.A1(\fmeasurment_nand4_ros.cycle_count[7] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0508_));
 sky130_fd_sc_hd__a221o_1 _1195_ (.A1(net321),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net334),
    .C1(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_4 _1196_ (.A(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0509_));
 sky130_fd_sc_hd__o221a_1 _1197_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[8] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[8] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0510_));
 sky130_fd_sc_hd__o211a_1 _1198_ (.A1(\fmeasurment_nand4_ros.cycle_count[8] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0511_));
 sky130_fd_sc_hd__a221o_1 _1199_ (.A1(\shift_register[8] ),
    .A2(_0509_),
    .B1(_0485_),
    .B2(net321),
    .C1(_0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_4 _1200_ (.A(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_4 _1201_ (.A(\ena_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0513_));
 sky130_fd_sc_hd__o221a_1 _1202_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[9] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[9] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0514_));
 sky130_fd_sc_hd__o211a_1 _1203_ (.A1(\fmeasurment_nand4_ros.cycle_count[9] ),
    .A2(_0487_),
    .B1(_0491_),
    .C1(_0514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0515_));
 sky130_fd_sc_hd__a221o_1 _1204_ (.A1(net332),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net335),
    .C1(_0515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__buf_2 _1205_ (.A(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_4 _1206_ (.A(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_4 _1207_ (.A(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0518_));
 sky130_fd_sc_hd__o221a_1 _1208_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[10] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[10] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0519_));
 sky130_fd_sc_hd__o211a_1 _1209_ (.A1(\fmeasurment_nand4_ros.cycle_count[10] ),
    .A2(_0487_),
    .B1(_0516_),
    .C1(_0519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0520_));
 sky130_fd_sc_hd__a221o_1 _1210_ (.A1(net326),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net332),
    .C1(_0520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_4 _1211_ (.A(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0521_));
 sky130_fd_sc_hd__o221a_1 _1212_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[11] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[11] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0522_));
 sky130_fd_sc_hd__o211a_1 _1213_ (.A1(\fmeasurment_nand4_ros.cycle_count[11] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0523_));
 sky130_fd_sc_hd__a221o_1 _1214_ (.A1(\shift_register[11] ),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net326),
    .C1(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__o221a_1 _1215_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[12] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[12] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0524_));
 sky130_fd_sc_hd__o211a_1 _1216_ (.A1(\fmeasurment_nand4_ros.cycle_count[12] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0525_));
 sky130_fd_sc_hd__a221o_1 _1217_ (.A1(\shift_register[12] ),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net336),
    .C1(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__o221a_1 _1218_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[13] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[13] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0526_));
 sky130_fd_sc_hd__o211a_1 _1219_ (.A1(\fmeasurment_nand4_ros.cycle_count[13] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0527_));
 sky130_fd_sc_hd__a221o_1 _1220_ (.A1(net328),
    .A2(_0509_),
    .B1(_0512_),
    .B2(\shift_register[12] ),
    .C1(_0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__o221a_1 _1221_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[14] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[14] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0528_));
 sky130_fd_sc_hd__o211a_1 _1222_ (.A1(\fmeasurment_nand4_ros.cycle_count[14] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0529_));
 sky130_fd_sc_hd__a221o_1 _1223_ (.A1(net339),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net328),
    .C1(_0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__o221a_1 _1224_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[15] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[15] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0530_));
 sky130_fd_sc_hd__o211a_1 _1225_ (.A1(\fmeasurment_nand4_ros.cycle_count[15] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0531_));
 sky130_fd_sc_hd__a221o_1 _1226_ (.A1(net323),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net339),
    .C1(_0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__o221a_1 _1227_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[16] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[16] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0532_));
 sky130_fd_sc_hd__o211a_1 _1228_ (.A1(\fmeasurment_nand4_ros.cycle_count[16] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0533_));
 sky130_fd_sc_hd__a221o_1 _1229_ (.A1(\shift_register[16] ),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net323),
    .C1(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__o221a_1 _1230_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[17] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[17] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0534_));
 sky130_fd_sc_hd__o211a_1 _1231_ (.A1(\fmeasurment_nand4_ros.cycle_count[17] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0535_));
 sky130_fd_sc_hd__a221o_1 _1232_ (.A1(\shift_register[17] ),
    .A2(_0509_),
    .B1(_0512_),
    .B2(net344),
    .C1(_0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__o221a_1 _1233_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[18] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[18] ),
    .C1(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0536_));
 sky130_fd_sc_hd__o211a_1 _1234_ (.A1(\fmeasurment_nand4_ros.cycle_count[18] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0537_));
 sky130_fd_sc_hd__a221o_1 _1235_ (.A1(net325),
    .A2(_0482_),
    .B1(_0512_),
    .B2(net347),
    .C1(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__o221a_1 _1236_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[19] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[19] ),
    .C1(\ena_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0538_));
 sky130_fd_sc_hd__o211a_1 _1237_ (.A1(\fmeasurment_nand4_ros.cycle_count[19] ),
    .A2(_0521_),
    .B1(_0516_),
    .C1(_0538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0539_));
 sky130_fd_sc_hd__a221o_1 _1238_ (.A1(net317),
    .A2(_0482_),
    .B1(_0484_),
    .B2(net325),
    .C1(_0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__and2_1 _1239_ (.A(_0494_),
    .B(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0540_));
 sky130_fd_sc_hd__a221o_1 _1240_ (.A1(\shift_register[21] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(net314),
    .C1(_0540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__a221o_1 _1241_ (.A1(\shift_register[23] ),
    .A2(_0482_),
    .B1(_0484_),
    .B2(net342),
    .C1(_0540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _1242_ (.A1(net314),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net317),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _1243_ (.A1(\shift_register[22] ),
    .A2(_0483_),
    .B1(_0485_),
    .B2(net319),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__o221a_1 _1244_ (.A1(\fmeasurment_einv_sub_ros.cycle_count[0] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(\fmeasurment_nand4_cap_ros.cycle_count[0] ),
    .C1(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0541_));
 sky130_fd_sc_hd__or2_1 _1245_ (.A(\fmeasurment_nand4_ros.cycle_count[0] ),
    .B(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0542_));
 sky130_fd_sc_hd__a32o_1 _1246_ (.A1(_0491_),
    .A2(_0541_),
    .A3(_0542_),
    .B1(_0483_),
    .B2(net316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__buf_4 _1247_ (.A(\ros_nand4.nets_notouch_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0543_));
 sky130_fd_sc_hd__buf_4 _1248_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0544_));
 sky130_fd_sc_hd__inv_2 _1249_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _1250_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1251_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1252_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1253_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1254_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1255_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1256_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1257_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1258_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_4 _1259_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0545_));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1261_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1262_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1263_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1264_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1266_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1267_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1268_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1269_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _1270_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0546_));
 sky130_fd_sc_hd__inv_2 _1271_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1272_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1273_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1274_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1275_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1276_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0025_));
 sky130_fd_sc_hd__buf_4 _1277_ (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0547_));
 sky130_fd_sc_hd__buf_4 _1278_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0548_));
 sky130_fd_sc_hd__inv_2 _1279_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1280_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1281_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1282_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1283_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1284_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1285_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1286_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1287_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0035_));
 sky130_fd_sc_hd__buf_4 _1289_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0549_));
 sky130_fd_sc_hd__inv_2 _1290_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1291_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1292_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1293_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1294_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1295_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1296_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1297_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1298_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1299_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1300_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1301_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1302_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0049_));
 sky130_fd_sc_hd__buf_4 _1304_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0550_));
 sky130_fd_sc_hd__inv_2 _1305_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1306_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1307_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1308_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1309_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1310_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1311_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1312_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1313_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1314_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1315_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1316_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1317_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1318_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1319_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1320_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0065_));
 sky130_fd_sc_hd__buf_4 _1321_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0551_));
 sky130_fd_sc_hd__inv_2 _1322_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1323_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1324_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1325_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1326_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1328_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1329_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1330_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1331_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0075_));
 sky130_fd_sc_hd__buf_4 _1332_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0552_));
 sky130_fd_sc_hd__inv_2 _1333_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1334_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1335_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1336_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1337_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1338_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1339_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1340_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1341_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1342_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1343_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1344_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1345_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1346_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1347_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1348_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0091_));
 sky130_fd_sc_hd__buf_4 _1349_ (.A(\ros_einv_sub.nets_notouch_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0553_));
 sky130_fd_sc_hd__buf_4 _1350_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0554_));
 sky130_fd_sc_hd__inv_2 _1351_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1352_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1353_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1354_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1355_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1359_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1360_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0101_));
 sky130_fd_sc_hd__buf_4 _1361_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0555_));
 sky130_fd_sc_hd__inv_2 _1362_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1363_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1364_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1365_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1366_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1367_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1368_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1369_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1370_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1371_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0111_));
 sky130_fd_sc_hd__buf_4 _1372_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0556_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1374_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1375_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1376_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1377_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1378_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1379_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1381_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1382_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0121_));
 sky130_fd_sc_hd__buf_4 _1383_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0557_));
 sky130_fd_sc_hd__inv_2 _1384_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1385_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1386_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1387_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1388_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1389_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1390_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1391_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1392_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1393_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1394_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1395_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1396_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1397_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1398_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1399_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0137_));
 sky130_fd_sc_hd__dfxtp_1 _1400_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1401_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1402_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1403_ (.CLK(clknet_2_3__leaf_clk),
    .D(net341),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1404_ (.CLK(clknet_2_3__leaf_clk),
    .D(net331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1405_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1406_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1407_ (.CLK(clknet_2_1__leaf_clk),
    .D(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1408_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1409_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1410_ (.CLK(clknet_2_1__leaf_clk),
    .D(net327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1411_ (.CLK(clknet_2_1__leaf_clk),
    .D(net337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1412_ (.CLK(clknet_2_1__leaf_clk),
    .D(net329),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1413_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1414_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1415_ (.CLK(clknet_2_0__leaf_clk),
    .D(net324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1416_ (.CLK(clknet_2_0__leaf_clk),
    .D(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1417_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1418_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1419_ (.CLK(clknet_2_2__leaf_clk),
    .D(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1420_ (.CLK(clknet_2_2__leaf_clk),
    .D(net343),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1421_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1422_ (.CLK(clknet_2_2__leaf_clk),
    .D(net320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1423_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\shift_register[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1424_ (.CLK(clknet_2_3__leaf_clk),
    .D(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\send_counter_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1425_ (.CLK(clknet_2_2__leaf_clk),
    .D(net311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\send_counter_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1426_ (.CLK(clknet_2_3__leaf_clk),
    .D(net312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\send_counter_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1427_ (.CLK(clknet_2_0__leaf_clk),
    .D(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ena_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1428_ (.CLK(clknet_2_0__leaf_clk),
    .D(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ena_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1429_ (.CLK(clknet_2_1__leaf_clk),
    .D(net310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ena_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1430_ (.CLK(_0000_),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.reset_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1431_ (.CLK(_0001_),
    .D(\fmeasurment_nand4_ros.reset_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.reset_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(_0002_),
    .D(\fmeasurment_nand4_ros.reset_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.reset_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(_0003_),
    .D(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1434_ (.CLK(_0004_),
    .D(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1435_ (.CLK(_0005_),
    .D(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1436_ (.CLK(_0006_),
    .D(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1437_ (.CLK(_0007_),
    .D(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1438_ (.CLK(_0008_),
    .D(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1439_ (.CLK(_0009_),
    .D(_0168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1440_ (.CLK(_0010_),
    .D(_0169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1441_ (.CLK(_0011_),
    .D(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1442_ (.CLK(_0012_),
    .D(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1443_ (.CLK(_0013_),
    .D(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1444_ (.CLK(_0014_),
    .D(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1445_ (.CLK(_0015_),
    .D(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1446_ (.CLK(_0016_),
    .D(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1447_ (.CLK(_0017_),
    .D(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1448_ (.CLK(_0018_),
    .D(_0177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1449_ (.CLK(_0019_),
    .D(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1450_ (.CLK(_0020_),
    .D(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(_0021_),
    .D(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(_0022_),
    .D(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.counts[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(_0023_),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.latch_counter_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1454_ (.CLK(_0024_),
    .D(\fmeasurment_nand4_ros.latch_counter_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.latch_counter_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1455_ (.CLK(_0025_),
    .D(\fmeasurment_nand4_ros.latch_counter_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.latch_counter_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1456_ (.CLK(_0026_),
    .D(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(_0027_),
    .D(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(_0028_),
    .D(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(_0029_),
    .D(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(_0030_),
    .D(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(_0031_),
    .D(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(_0032_),
    .D(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(_0033_),
    .D(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(_0034_),
    .D(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(_0035_),
    .D(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(_0036_),
    .D(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(_0037_),
    .D(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1468_ (.CLK(_0038_),
    .D(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1469_ (.CLK(_0039_),
    .D(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1470_ (.CLK(_0040_),
    .D(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1471_ (.CLK(_0041_),
    .D(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1472_ (.CLK(_0042_),
    .D(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1473_ (.CLK(_0043_),
    .D(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1474_ (.CLK(_0044_),
    .D(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1475_ (.CLK(_0045_),
    .D(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.cycle_count[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1476_ (.CLK(_0046_),
    .D(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1477_ (.CLK(_0047_),
    .D(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1478_ (.CLK(_0048_),
    .D(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1479_ (.CLK(_0049_),
    .D(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1480_ (.CLK(_0050_),
    .D(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1481_ (.CLK(_0051_),
    .D(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1482_ (.CLK(_0052_),
    .D(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1483_ (.CLK(_0053_),
    .D(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1484_ (.CLK(_0054_),
    .D(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1485_ (.CLK(_0055_),
    .D(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1486_ (.CLK(_0056_),
    .D(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1487_ (.CLK(_0057_),
    .D(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1488_ (.CLK(_0058_),
    .D(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1489_ (.CLK(_0059_),
    .D(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1490_ (.CLK(_0060_),
    .D(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1491_ (.CLK(_0061_),
    .D(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1492_ (.CLK(_0062_),
    .D(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1493_ (.CLK(_0063_),
    .D(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1494_ (.CLK(_0064_),
    .D(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1495_ (.CLK(_0065_),
    .D(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_ros.cycle_count[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1496_ (.CLK(_0066_),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.reset_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1497_ (.CLK(_0067_),
    .D(\fmeasurment_nand4_cap_ros.reset_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.reset_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1498_ (.CLK(_0068_),
    .D(\fmeasurment_nand4_cap_ros.reset_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.reset_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1499_ (.CLK(_0069_),
    .D(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1500_ (.CLK(_0070_),
    .D(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1501_ (.CLK(_0071_),
    .D(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1502_ (.CLK(_0072_),
    .D(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1503_ (.CLK(_0073_),
    .D(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1504_ (.CLK(_0074_),
    .D(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1505_ (.CLK(_0075_),
    .D(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1506_ (.CLK(_0076_),
    .D(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1507_ (.CLK(_0077_),
    .D(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1508_ (.CLK(_0078_),
    .D(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1509_ (.CLK(_0079_),
    .D(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1510_ (.CLK(_0080_),
    .D(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1511_ (.CLK(_0081_),
    .D(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1512_ (.CLK(_0082_),
    .D(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1513_ (.CLK(_0083_),
    .D(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1514_ (.CLK(_0084_),
    .D(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1515_ (.CLK(_0085_),
    .D(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1516_ (.CLK(_0086_),
    .D(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1517_ (.CLK(_0087_),
    .D(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1518_ (.CLK(_0088_),
    .D(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.counts[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1519_ (.CLK(_0089_),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.latch_counter_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1520_ (.CLK(_0090_),
    .D(\fmeasurment_nand4_cap_ros.latch_counter_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.latch_counter_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1521_ (.CLK(_0091_),
    .D(\fmeasurment_nand4_cap_ros.latch_counter_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_nand4_cap_ros.latch_counter_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1522_ (.CLK(_0092_),
    .D(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1523_ (.CLK(_0093_),
    .D(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1524_ (.CLK(_0094_),
    .D(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1525_ (.CLK(_0095_),
    .D(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1526_ (.CLK(_0096_),
    .D(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1527_ (.CLK(_0097_),
    .D(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1528_ (.CLK(_0098_),
    .D(_0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1529_ (.CLK(_0099_),
    .D(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1530_ (.CLK(_0100_),
    .D(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1531_ (.CLK(_0101_),
    .D(_0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1532_ (.CLK(_0102_),
    .D(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1533_ (.CLK(_0103_),
    .D(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1534_ (.CLK(_0104_),
    .D(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1535_ (.CLK(_0105_),
    .D(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1536_ (.CLK(_0106_),
    .D(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1537_ (.CLK(_0107_),
    .D(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1538_ (.CLK(_0108_),
    .D(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1539_ (.CLK(_0109_),
    .D(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1540_ (.CLK(_0110_),
    .D(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1541_ (.CLK(_0111_),
    .D(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.cycle_count[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1542_ (.CLK(_0112_),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.reset_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1543_ (.CLK(_0113_),
    .D(\fmeasurment_einv_sub_ros.reset_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.reset_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1544_ (.CLK(_0114_),
    .D(\fmeasurment_einv_sub_ros.reset_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.reset_syncs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1545_ (.CLK(_0115_),
    .D(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1546_ (.CLK(_0116_),
    .D(_0263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1547_ (.CLK(_0117_),
    .D(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1548_ (.CLK(_0118_),
    .D(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1549_ (.CLK(_0119_),
    .D(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1550_ (.CLK(_0120_),
    .D(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1551_ (.CLK(_0121_),
    .D(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1552_ (.CLK(_0122_),
    .D(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1553_ (.CLK(_0123_),
    .D(_0270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1554_ (.CLK(_0124_),
    .D(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1555_ (.CLK(_0125_),
    .D(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1556_ (.CLK(_0126_),
    .D(_0273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1557_ (.CLK(_0127_),
    .D(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1558_ (.CLK(_0128_),
    .D(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1559_ (.CLK(_0129_),
    .D(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1560_ (.CLK(_0130_),
    .D(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1561_ (.CLK(_0131_),
    .D(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1562_ (.CLK(_0132_),
    .D(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1563_ (.CLK(_0133_),
    .D(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1564_ (.CLK(_0134_),
    .D(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.counts[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1565_ (.CLK(_0135_),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.latch_counter_syncs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1566_ (.CLK(_0136_),
    .D(\fmeasurment_einv_sub_ros.latch_counter_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.latch_counter_syncs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1567_ (.CLK(_0137_),
    .D(\fmeasurment_einv_sub_ros.latch_counter_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fmeasurment_einv_sub_ros.latch_counter_syncs[2] ));
 sky130_fd_sc_hd__buf_2 _1868_ (.A(data_stream),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _1869_ (.A(\fmeasurment_einv_sub_ros.divided_clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _1870_ (.A(\fmeasurment_nand4_cap_ros.divided_clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _1871_ (.A(\fmeasurment_nand4_ros.divided_clk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\ena_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\shift_register[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\shift_register[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\shift_register[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\shift_register[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\shift_register[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\shift_register[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\send_counter_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\shift_register[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\shift_register[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\shift_register[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\shift_register[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\shift_register[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\shift_register[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ena_syncs[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\send_counter_syncs[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\shift_register[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\shift_register[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\shift_register[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\shift_register[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\shift_register[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\shift_register[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\ena_syncs[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\shift_register[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\shift_register[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\shift_register[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\shift_register[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__nand2_1 \ros_einv_sub.fstage  (.A(\ros_einv_sub.nets_notouch_[24] ),
    .B(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[0] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[0].genblk1[0].tristage  (.A(\ros_einv_sub.nets_notouch_[0] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[1] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[0].genblk1[1].tristage  (.A(\ros_einv_sub.nets_notouch_[1] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[2] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[0].genblk1[2].tristage  (.A(\ros_einv_sub.nets_notouch_[2] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[3] ));
 sky130_fd_sc_hd__inv_1 \ros_einv_sub.genblk1[0].stage  (.A(\ros_einv_sub.nets_notouch_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[4] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[1].genblk1[0].tristage  (.A(\ros_einv_sub.nets_notouch_[4] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[5] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[1].genblk1[1].tristage  (.A(\ros_einv_sub.nets_notouch_[5] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[6] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[1].genblk1[2].tristage  (.A(\ros_einv_sub.nets_notouch_[6] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[7] ));
 sky130_fd_sc_hd__inv_1 \ros_einv_sub.genblk1[1].stage  (.A(\ros_einv_sub.nets_notouch_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[8] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[2].genblk1[0].tristage  (.A(\ros_einv_sub.nets_notouch_[8] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[9] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[2].genblk1[1].tristage  (.A(\ros_einv_sub.nets_notouch_[9] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[10] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[2].genblk1[2].tristage  (.A(\ros_einv_sub.nets_notouch_[10] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[11] ));
 sky130_fd_sc_hd__inv_1 \ros_einv_sub.genblk1[2].stage  (.A(\ros_einv_sub.nets_notouch_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[12] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[3].genblk1[0].tristage  (.A(\ros_einv_sub.nets_notouch_[12] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[13] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[3].genblk1[1].tristage  (.A(\ros_einv_sub.nets_notouch_[13] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[14] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[3].genblk1[2].tristage  (.A(\ros_einv_sub.nets_notouch_[14] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[15] ));
 sky130_fd_sc_hd__inv_1 \ros_einv_sub.genblk1[3].stage  (.A(\ros_einv_sub.nets_notouch_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[16] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[4].genblk1[0].tristage  (.A(\ros_einv_sub.nets_notouch_[16] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[17] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[4].genblk1[1].tristage  (.A(\ros_einv_sub.nets_notouch_[17] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[18] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[4].genblk1[2].tristage  (.A(\ros_einv_sub.nets_notouch_[18] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[19] ));
 sky130_fd_sc_hd__inv_1 \ros_einv_sub.genblk1[4].stage  (.A(\ros_einv_sub.nets_notouch_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[20] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[5].genblk1[0].tristage  (.A(\ros_einv_sub.nets_notouch_[20] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[21] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[5].genblk1[1].tristage  (.A(\ros_einv_sub.nets_notouch_[21] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[22] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.genblk1[5].genblk1[2].tristage  (.A(\ros_einv_sub.nets_notouch_[22] ),
    .TE(\ros_einv_sub.sub_voltage_notouch_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.nets_notouch_[23] ));
 sky130_fd_sc_hd__inv_1 \ros_einv_sub.genblk1[5].stage  (.A(\ros_einv_sub.nets_notouch_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_einv_sub.nets_notouch_[24] ));
 sky130_fd_sc_hd__einvp_1 \ros_einv_sub.sub_generator  (.A(\ros_einv_sub.sub_voltage_notouch_ ),
    .TE(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\ros_einv_sub.sub_voltage_notouch_ ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.fstage  (.A(net1),
    .B(\ros_nand4.nets_notouch_[66] ),
    .C(\ros_nand4.nets_notouch_[66] ),
    .D(\ros_nand4.nets_notouch_[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[0] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[10].stage  (.A(\ros_nand4.nets_notouch_[9] ),
    .B(\ros_nand4.nets_notouch_[9] ),
    .C(\ros_nand4.nets_notouch_[9] ),
    .D(\ros_nand4.nets_notouch_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[10] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[11].stage  (.A(\ros_nand4.nets_notouch_[10] ),
    .B(\ros_nand4.nets_notouch_[10] ),
    .C(\ros_nand4.nets_notouch_[10] ),
    .D(\ros_nand4.nets_notouch_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[11] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[12].stage  (.A(\ros_nand4.nets_notouch_[11] ),
    .B(\ros_nand4.nets_notouch_[11] ),
    .C(\ros_nand4.nets_notouch_[11] ),
    .D(\ros_nand4.nets_notouch_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[12] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[13].stage  (.A(\ros_nand4.nets_notouch_[12] ),
    .B(\ros_nand4.nets_notouch_[12] ),
    .C(\ros_nand4.nets_notouch_[12] ),
    .D(\ros_nand4.nets_notouch_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[13] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[14].stage  (.A(\ros_nand4.nets_notouch_[13] ),
    .B(\ros_nand4.nets_notouch_[13] ),
    .C(\ros_nand4.nets_notouch_[13] ),
    .D(\ros_nand4.nets_notouch_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[14] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[15].stage  (.A(\ros_nand4.nets_notouch_[14] ),
    .B(\ros_nand4.nets_notouch_[14] ),
    .C(\ros_nand4.nets_notouch_[14] ),
    .D(\ros_nand4.nets_notouch_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[15] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[16].stage  (.A(\ros_nand4.nets_notouch_[15] ),
    .B(\ros_nand4.nets_notouch_[15] ),
    .C(\ros_nand4.nets_notouch_[15] ),
    .D(\ros_nand4.nets_notouch_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[16] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[17].stage  (.A(\ros_nand4.nets_notouch_[16] ),
    .B(\ros_nand4.nets_notouch_[16] ),
    .C(\ros_nand4.nets_notouch_[16] ),
    .D(\ros_nand4.nets_notouch_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[17] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[18].stage  (.A(\ros_nand4.nets_notouch_[17] ),
    .B(\ros_nand4.nets_notouch_[17] ),
    .C(\ros_nand4.nets_notouch_[17] ),
    .D(\ros_nand4.nets_notouch_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[18] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[19].stage  (.A(\ros_nand4.nets_notouch_[18] ),
    .B(\ros_nand4.nets_notouch_[18] ),
    .C(\ros_nand4.nets_notouch_[18] ),
    .D(\ros_nand4.nets_notouch_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[19] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[1].stage  (.A(\ros_nand4.nets_notouch_[0] ),
    .B(\ros_nand4.nets_notouch_[0] ),
    .C(\ros_nand4.nets_notouch_[0] ),
    .D(\ros_nand4.nets_notouch_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[1] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[20].stage  (.A(\ros_nand4.nets_notouch_[19] ),
    .B(\ros_nand4.nets_notouch_[19] ),
    .C(\ros_nand4.nets_notouch_[19] ),
    .D(\ros_nand4.nets_notouch_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[20] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[21].stage  (.A(\ros_nand4.nets_notouch_[20] ),
    .B(\ros_nand4.nets_notouch_[20] ),
    .C(\ros_nand4.nets_notouch_[20] ),
    .D(\ros_nand4.nets_notouch_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[21] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[22].stage  (.A(\ros_nand4.nets_notouch_[21] ),
    .B(\ros_nand4.nets_notouch_[21] ),
    .C(\ros_nand4.nets_notouch_[21] ),
    .D(\ros_nand4.nets_notouch_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[22] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[23].stage  (.A(\ros_nand4.nets_notouch_[22] ),
    .B(\ros_nand4.nets_notouch_[22] ),
    .C(\ros_nand4.nets_notouch_[22] ),
    .D(\ros_nand4.nets_notouch_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[23] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[24].stage  (.A(\ros_nand4.nets_notouch_[23] ),
    .B(\ros_nand4.nets_notouch_[23] ),
    .C(\ros_nand4.nets_notouch_[23] ),
    .D(\ros_nand4.nets_notouch_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[24] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[25].stage  (.A(\ros_nand4.nets_notouch_[24] ),
    .B(\ros_nand4.nets_notouch_[24] ),
    .C(\ros_nand4.nets_notouch_[24] ),
    .D(\ros_nand4.nets_notouch_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[25] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[26].stage  (.A(\ros_nand4.nets_notouch_[25] ),
    .B(\ros_nand4.nets_notouch_[25] ),
    .C(\ros_nand4.nets_notouch_[25] ),
    .D(\ros_nand4.nets_notouch_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[26] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[27].stage  (.A(\ros_nand4.nets_notouch_[26] ),
    .B(\ros_nand4.nets_notouch_[26] ),
    .C(\ros_nand4.nets_notouch_[26] ),
    .D(\ros_nand4.nets_notouch_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[27] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[28].stage  (.A(\ros_nand4.nets_notouch_[27] ),
    .B(\ros_nand4.nets_notouch_[27] ),
    .C(\ros_nand4.nets_notouch_[27] ),
    .D(\ros_nand4.nets_notouch_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[28] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[29].stage  (.A(\ros_nand4.nets_notouch_[28] ),
    .B(\ros_nand4.nets_notouch_[28] ),
    .C(\ros_nand4.nets_notouch_[28] ),
    .D(\ros_nand4.nets_notouch_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[29] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[2].stage  (.A(\ros_nand4.nets_notouch_[1] ),
    .B(\ros_nand4.nets_notouch_[1] ),
    .C(\ros_nand4.nets_notouch_[1] ),
    .D(\ros_nand4.nets_notouch_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[2] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[30].stage  (.A(\ros_nand4.nets_notouch_[29] ),
    .B(\ros_nand4.nets_notouch_[29] ),
    .C(\ros_nand4.nets_notouch_[29] ),
    .D(\ros_nand4.nets_notouch_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[30] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[31].stage  (.A(\ros_nand4.nets_notouch_[30] ),
    .B(\ros_nand4.nets_notouch_[30] ),
    .C(\ros_nand4.nets_notouch_[30] ),
    .D(\ros_nand4.nets_notouch_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[31] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[32].stage  (.A(\ros_nand4.nets_notouch_[31] ),
    .B(\ros_nand4.nets_notouch_[31] ),
    .C(\ros_nand4.nets_notouch_[31] ),
    .D(\ros_nand4.nets_notouch_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[32] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[33].stage  (.A(\ros_nand4.nets_notouch_[32] ),
    .B(\ros_nand4.nets_notouch_[32] ),
    .C(\ros_nand4.nets_notouch_[32] ),
    .D(\ros_nand4.nets_notouch_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[33] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[34].stage  (.A(\ros_nand4.nets_notouch_[33] ),
    .B(\ros_nand4.nets_notouch_[33] ),
    .C(\ros_nand4.nets_notouch_[33] ),
    .D(\ros_nand4.nets_notouch_[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[34] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[35].stage  (.A(\ros_nand4.nets_notouch_[34] ),
    .B(\ros_nand4.nets_notouch_[34] ),
    .C(\ros_nand4.nets_notouch_[34] ),
    .D(\ros_nand4.nets_notouch_[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[35] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[36].stage  (.A(\ros_nand4.nets_notouch_[35] ),
    .B(\ros_nand4.nets_notouch_[35] ),
    .C(\ros_nand4.nets_notouch_[35] ),
    .D(\ros_nand4.nets_notouch_[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[36] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[37].stage  (.A(\ros_nand4.nets_notouch_[36] ),
    .B(\ros_nand4.nets_notouch_[36] ),
    .C(\ros_nand4.nets_notouch_[36] ),
    .D(\ros_nand4.nets_notouch_[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[37] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[38].stage  (.A(\ros_nand4.nets_notouch_[37] ),
    .B(\ros_nand4.nets_notouch_[37] ),
    .C(\ros_nand4.nets_notouch_[37] ),
    .D(\ros_nand4.nets_notouch_[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[38] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[39].stage  (.A(\ros_nand4.nets_notouch_[38] ),
    .B(\ros_nand4.nets_notouch_[38] ),
    .C(\ros_nand4.nets_notouch_[38] ),
    .D(\ros_nand4.nets_notouch_[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[39] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[3].stage  (.A(\ros_nand4.nets_notouch_[2] ),
    .B(\ros_nand4.nets_notouch_[2] ),
    .C(\ros_nand4.nets_notouch_[2] ),
    .D(\ros_nand4.nets_notouch_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[3] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[40].stage  (.A(\ros_nand4.nets_notouch_[39] ),
    .B(\ros_nand4.nets_notouch_[39] ),
    .C(\ros_nand4.nets_notouch_[39] ),
    .D(\ros_nand4.nets_notouch_[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[40] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[41].stage  (.A(\ros_nand4.nets_notouch_[40] ),
    .B(\ros_nand4.nets_notouch_[40] ),
    .C(\ros_nand4.nets_notouch_[40] ),
    .D(\ros_nand4.nets_notouch_[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[41] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[42].stage  (.A(\ros_nand4.nets_notouch_[41] ),
    .B(\ros_nand4.nets_notouch_[41] ),
    .C(\ros_nand4.nets_notouch_[41] ),
    .D(\ros_nand4.nets_notouch_[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[42] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[43].stage  (.A(\ros_nand4.nets_notouch_[42] ),
    .B(\ros_nand4.nets_notouch_[42] ),
    .C(\ros_nand4.nets_notouch_[42] ),
    .D(\ros_nand4.nets_notouch_[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[43] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[44].stage  (.A(\ros_nand4.nets_notouch_[43] ),
    .B(\ros_nand4.nets_notouch_[43] ),
    .C(\ros_nand4.nets_notouch_[43] ),
    .D(\ros_nand4.nets_notouch_[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[44] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[45].stage  (.A(\ros_nand4.nets_notouch_[44] ),
    .B(\ros_nand4.nets_notouch_[44] ),
    .C(\ros_nand4.nets_notouch_[44] ),
    .D(\ros_nand4.nets_notouch_[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[45] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[46].stage  (.A(\ros_nand4.nets_notouch_[45] ),
    .B(\ros_nand4.nets_notouch_[45] ),
    .C(\ros_nand4.nets_notouch_[45] ),
    .D(\ros_nand4.nets_notouch_[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[46] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[47].stage  (.A(\ros_nand4.nets_notouch_[46] ),
    .B(\ros_nand4.nets_notouch_[46] ),
    .C(\ros_nand4.nets_notouch_[46] ),
    .D(\ros_nand4.nets_notouch_[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[47] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[48].stage  (.A(\ros_nand4.nets_notouch_[47] ),
    .B(\ros_nand4.nets_notouch_[47] ),
    .C(\ros_nand4.nets_notouch_[47] ),
    .D(\ros_nand4.nets_notouch_[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[48] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[49].stage  (.A(\ros_nand4.nets_notouch_[48] ),
    .B(\ros_nand4.nets_notouch_[48] ),
    .C(\ros_nand4.nets_notouch_[48] ),
    .D(\ros_nand4.nets_notouch_[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[49] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[4].stage  (.A(\ros_nand4.nets_notouch_[3] ),
    .B(\ros_nand4.nets_notouch_[3] ),
    .C(\ros_nand4.nets_notouch_[3] ),
    .D(\ros_nand4.nets_notouch_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[4] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[50].stage  (.A(\ros_nand4.nets_notouch_[49] ),
    .B(\ros_nand4.nets_notouch_[49] ),
    .C(\ros_nand4.nets_notouch_[49] ),
    .D(\ros_nand4.nets_notouch_[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[50] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[51].stage  (.A(\ros_nand4.nets_notouch_[50] ),
    .B(\ros_nand4.nets_notouch_[50] ),
    .C(\ros_nand4.nets_notouch_[50] ),
    .D(\ros_nand4.nets_notouch_[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[51] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[52].stage  (.A(\ros_nand4.nets_notouch_[51] ),
    .B(\ros_nand4.nets_notouch_[51] ),
    .C(\ros_nand4.nets_notouch_[51] ),
    .D(\ros_nand4.nets_notouch_[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[52] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[53].stage  (.A(\ros_nand4.nets_notouch_[52] ),
    .B(\ros_nand4.nets_notouch_[52] ),
    .C(\ros_nand4.nets_notouch_[52] ),
    .D(\ros_nand4.nets_notouch_[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[53] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[54].stage  (.A(\ros_nand4.nets_notouch_[53] ),
    .B(\ros_nand4.nets_notouch_[53] ),
    .C(\ros_nand4.nets_notouch_[53] ),
    .D(\ros_nand4.nets_notouch_[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[54] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[55].stage  (.A(\ros_nand4.nets_notouch_[54] ),
    .B(\ros_nand4.nets_notouch_[54] ),
    .C(\ros_nand4.nets_notouch_[54] ),
    .D(\ros_nand4.nets_notouch_[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[55] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[56].stage  (.A(\ros_nand4.nets_notouch_[55] ),
    .B(\ros_nand4.nets_notouch_[55] ),
    .C(\ros_nand4.nets_notouch_[55] ),
    .D(\ros_nand4.nets_notouch_[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[56] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[57].stage  (.A(\ros_nand4.nets_notouch_[56] ),
    .B(\ros_nand4.nets_notouch_[56] ),
    .C(\ros_nand4.nets_notouch_[56] ),
    .D(\ros_nand4.nets_notouch_[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[57] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[58].stage  (.A(\ros_nand4.nets_notouch_[57] ),
    .B(\ros_nand4.nets_notouch_[57] ),
    .C(\ros_nand4.nets_notouch_[57] ),
    .D(\ros_nand4.nets_notouch_[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[58] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[59].stage  (.A(\ros_nand4.nets_notouch_[58] ),
    .B(\ros_nand4.nets_notouch_[58] ),
    .C(\ros_nand4.nets_notouch_[58] ),
    .D(\ros_nand4.nets_notouch_[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[59] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[5].stage  (.A(\ros_nand4.nets_notouch_[4] ),
    .B(\ros_nand4.nets_notouch_[4] ),
    .C(\ros_nand4.nets_notouch_[4] ),
    .D(\ros_nand4.nets_notouch_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[5] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[60].stage  (.A(\ros_nand4.nets_notouch_[59] ),
    .B(\ros_nand4.nets_notouch_[59] ),
    .C(\ros_nand4.nets_notouch_[59] ),
    .D(\ros_nand4.nets_notouch_[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[60] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[61].stage  (.A(\ros_nand4.nets_notouch_[60] ),
    .B(\ros_nand4.nets_notouch_[60] ),
    .C(\ros_nand4.nets_notouch_[60] ),
    .D(\ros_nand4.nets_notouch_[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[61] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[62].stage  (.A(\ros_nand4.nets_notouch_[61] ),
    .B(\ros_nand4.nets_notouch_[61] ),
    .C(\ros_nand4.nets_notouch_[61] ),
    .D(\ros_nand4.nets_notouch_[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[62] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[63].stage  (.A(\ros_nand4.nets_notouch_[62] ),
    .B(\ros_nand4.nets_notouch_[62] ),
    .C(\ros_nand4.nets_notouch_[62] ),
    .D(\ros_nand4.nets_notouch_[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[63] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[64].stage  (.A(\ros_nand4.nets_notouch_[63] ),
    .B(\ros_nand4.nets_notouch_[63] ),
    .C(\ros_nand4.nets_notouch_[63] ),
    .D(\ros_nand4.nets_notouch_[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[64] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[65].stage  (.A(\ros_nand4.nets_notouch_[64] ),
    .B(\ros_nand4.nets_notouch_[64] ),
    .C(\ros_nand4.nets_notouch_[64] ),
    .D(\ros_nand4.nets_notouch_[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[65] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[66].stage  (.A(\ros_nand4.nets_notouch_[65] ),
    .B(\ros_nand4.nets_notouch_[65] ),
    .C(\ros_nand4.nets_notouch_[65] ),
    .D(\ros_nand4.nets_notouch_[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[66] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[6].stage  (.A(\ros_nand4.nets_notouch_[5] ),
    .B(\ros_nand4.nets_notouch_[5] ),
    .C(\ros_nand4.nets_notouch_[5] ),
    .D(\ros_nand4.nets_notouch_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[6] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[7].stage  (.A(\ros_nand4.nets_notouch_[6] ),
    .B(\ros_nand4.nets_notouch_[6] ),
    .C(\ros_nand4.nets_notouch_[6] ),
    .D(\ros_nand4.nets_notouch_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[7] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[8].stage  (.A(\ros_nand4.nets_notouch_[7] ),
    .B(\ros_nand4.nets_notouch_[7] ),
    .C(\ros_nand4.nets_notouch_[7] ),
    .D(\ros_nand4.nets_notouch_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[8] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4.genblk1[9].stage  (.A(\ros_nand4.nets_notouch_[8] ),
    .B(\ros_nand4.nets_notouch_[8] ),
    .C(\ros_nand4.nets_notouch_[8] ),
    .D(\ros_nand4.nets_notouch_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4.nets_notouch_[9] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.fstage  (.A(net1),
    .B(\ros_nand4_cap.nets_notouch_[34] ),
    .C(\ros_nand4_cap.nets_notouch_[34] ),
    .D(\ros_nand4_cap.nets_notouch_[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[0] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[10].stage  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(\ros_nand4_cap.nets_notouch_[9] ),
    .C(\ros_nand4_cap.nets_notouch_[9] ),
    .D(\ros_nand4_cap.nets_notouch_[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[10] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[11].stage  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(\ros_nand4_cap.nets_notouch_[10] ),
    .C(\ros_nand4_cap.nets_notouch_[10] ),
    .D(\ros_nand4_cap.nets_notouch_[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[11] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[12].stage  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(\ros_nand4_cap.nets_notouch_[11] ),
    .C(\ros_nand4_cap.nets_notouch_[11] ),
    .D(\ros_nand4_cap.nets_notouch_[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[12] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[13].stage  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(\ros_nand4_cap.nets_notouch_[12] ),
    .C(\ros_nand4_cap.nets_notouch_[12] ),
    .D(\ros_nand4_cap.nets_notouch_[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[13] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[14].stage  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(\ros_nand4_cap.nets_notouch_[13] ),
    .C(\ros_nand4_cap.nets_notouch_[13] ),
    .D(\ros_nand4_cap.nets_notouch_[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[14] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[15].stage  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(\ros_nand4_cap.nets_notouch_[14] ),
    .C(\ros_nand4_cap.nets_notouch_[14] ),
    .D(\ros_nand4_cap.nets_notouch_[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[15] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[16].stage  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(\ros_nand4_cap.nets_notouch_[15] ),
    .C(\ros_nand4_cap.nets_notouch_[15] ),
    .D(\ros_nand4_cap.nets_notouch_[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[16] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[17].stage  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(\ros_nand4_cap.nets_notouch_[16] ),
    .C(\ros_nand4_cap.nets_notouch_[16] ),
    .D(\ros_nand4_cap.nets_notouch_[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[17] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[18].stage  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(\ros_nand4_cap.nets_notouch_[17] ),
    .C(\ros_nand4_cap.nets_notouch_[17] ),
    .D(\ros_nand4_cap.nets_notouch_[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[18] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[19].stage  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(\ros_nand4_cap.nets_notouch_[18] ),
    .C(\ros_nand4_cap.nets_notouch_[18] ),
    .D(\ros_nand4_cap.nets_notouch_[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[19] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[1].stage  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(\ros_nand4_cap.nets_notouch_[0] ),
    .C(\ros_nand4_cap.nets_notouch_[0] ),
    .D(\ros_nand4_cap.nets_notouch_[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[1] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[20].stage  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(\ros_nand4_cap.nets_notouch_[19] ),
    .C(\ros_nand4_cap.nets_notouch_[19] ),
    .D(\ros_nand4_cap.nets_notouch_[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[20] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[21].stage  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(\ros_nand4_cap.nets_notouch_[20] ),
    .C(\ros_nand4_cap.nets_notouch_[20] ),
    .D(\ros_nand4_cap.nets_notouch_[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[21] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[22].stage  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(\ros_nand4_cap.nets_notouch_[21] ),
    .C(\ros_nand4_cap.nets_notouch_[21] ),
    .D(\ros_nand4_cap.nets_notouch_[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[22] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[23].stage  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(\ros_nand4_cap.nets_notouch_[22] ),
    .C(\ros_nand4_cap.nets_notouch_[22] ),
    .D(\ros_nand4_cap.nets_notouch_[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[23] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[24].stage  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(\ros_nand4_cap.nets_notouch_[23] ),
    .C(\ros_nand4_cap.nets_notouch_[23] ),
    .D(\ros_nand4_cap.nets_notouch_[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[24] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[25].stage  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(\ros_nand4_cap.nets_notouch_[24] ),
    .C(\ros_nand4_cap.nets_notouch_[24] ),
    .D(\ros_nand4_cap.nets_notouch_[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[25] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[26].stage  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(\ros_nand4_cap.nets_notouch_[25] ),
    .C(\ros_nand4_cap.nets_notouch_[25] ),
    .D(\ros_nand4_cap.nets_notouch_[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[26] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[27].stage  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(\ros_nand4_cap.nets_notouch_[26] ),
    .C(\ros_nand4_cap.nets_notouch_[26] ),
    .D(\ros_nand4_cap.nets_notouch_[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[27] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[28].stage  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(\ros_nand4_cap.nets_notouch_[27] ),
    .C(\ros_nand4_cap.nets_notouch_[27] ),
    .D(\ros_nand4_cap.nets_notouch_[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[28] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[29].stage  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(\ros_nand4_cap.nets_notouch_[28] ),
    .C(\ros_nand4_cap.nets_notouch_[28] ),
    .D(\ros_nand4_cap.nets_notouch_[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[29] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[2].stage  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(\ros_nand4_cap.nets_notouch_[1] ),
    .C(\ros_nand4_cap.nets_notouch_[1] ),
    .D(\ros_nand4_cap.nets_notouch_[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[2] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[30].stage  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(\ros_nand4_cap.nets_notouch_[29] ),
    .C(\ros_nand4_cap.nets_notouch_[29] ),
    .D(\ros_nand4_cap.nets_notouch_[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[30] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[31].stage  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(\ros_nand4_cap.nets_notouch_[30] ),
    .C(\ros_nand4_cap.nets_notouch_[30] ),
    .D(\ros_nand4_cap.nets_notouch_[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[31] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[32].stage  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(\ros_nand4_cap.nets_notouch_[31] ),
    .C(\ros_nand4_cap.nets_notouch_[31] ),
    .D(\ros_nand4_cap.nets_notouch_[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[32] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[33].stage  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(\ros_nand4_cap.nets_notouch_[32] ),
    .C(\ros_nand4_cap.nets_notouch_[32] ),
    .D(\ros_nand4_cap.nets_notouch_[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[33] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[34].stage  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(\ros_nand4_cap.nets_notouch_[33] ),
    .C(\ros_nand4_cap.nets_notouch_[33] ),
    .D(\ros_nand4_cap.nets_notouch_[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[34] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[3].stage  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(\ros_nand4_cap.nets_notouch_[2] ),
    .C(\ros_nand4_cap.nets_notouch_[2] ),
    .D(\ros_nand4_cap.nets_notouch_[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[3] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[4].stage  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(\ros_nand4_cap.nets_notouch_[3] ),
    .C(\ros_nand4_cap.nets_notouch_[3] ),
    .D(\ros_nand4_cap.nets_notouch_[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[4] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[5].stage  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(\ros_nand4_cap.nets_notouch_[4] ),
    .C(\ros_nand4_cap.nets_notouch_[4] ),
    .D(\ros_nand4_cap.nets_notouch_[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[5] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[6].stage  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(\ros_nand4_cap.nets_notouch_[5] ),
    .C(\ros_nand4_cap.nets_notouch_[5] ),
    .D(\ros_nand4_cap.nets_notouch_[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[6] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[7].stage  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(\ros_nand4_cap.nets_notouch_[6] ),
    .C(\ros_nand4_cap.nets_notouch_[6] ),
    .D(\ros_nand4_cap.nets_notouch_[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[7] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[8].stage  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(\ros_nand4_cap.nets_notouch_[7] ),
    .C(\ros_nand4_cap.nets_notouch_[7] ),
    .D(\ros_nand4_cap.nets_notouch_[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[8] ));
 sky130_fd_sc_hd__nand4_1 \ros_nand4_cap.genblk1[9].stage  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(\ros_nand4_cap.nets_notouch_[8] ),
    .C(\ros_nand4_cap.nets_notouch_[8] ),
    .D(\ros_nand4_cap.nets_notouch_[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.nets_notouch_[9] ));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[0] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[0].cap_10  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net10));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[1] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[1].cap_11  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net11));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[2] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[2].cap_12  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net12));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[3] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[3].cap_13  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net13));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[4] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[4].cap_14  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net14));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[5] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[5].cap_15  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net15));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[6] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[6].cap_16  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net16));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[0].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[0] ),
    .B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[7] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[0].genblk1[7].cap_17  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net17));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[80] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[0].cap_18  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net18));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[81] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[1].cap_19  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net19));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[82] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[2].cap_20  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net20));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[83] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[3].cap_21  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net21));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[84] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[4].cap_22  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net22));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[85] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[5].cap_23  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net23));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[86] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[6].cap_24  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net24));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[10].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[10] ),
    .B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[87] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[10].genblk1[7].cap_25  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net25));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[88] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[0].cap_26  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net26));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[89] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[1].cap_27  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net27));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[90] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[2].cap_28  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net28));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[91] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[3].cap_29  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net29));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[92] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[4].cap_30  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[93] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[5].cap_31  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[94] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[6].cap_32  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[11].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[11] ),
    .B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[95] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[11].genblk1[7].cap_33  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net33));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[96] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[0].cap_34  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net34));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[97] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[1].cap_35  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net35));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[98] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[2].cap_36  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net36));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[99] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[3].cap_37  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net37));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[100] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[4].cap_38  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net38));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[101] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[5].cap_39  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net39));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[102] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[6].cap_40  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net40));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[12].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[12] ),
    .B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[103] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[12].genblk1[7].cap_41  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net41));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[104] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[0].cap_42  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net42));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[105] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[1].cap_43  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net43));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[106] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[2].cap_44  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net44));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[107] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[3].cap_45  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net45));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[108] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[4].cap_46  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net46));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[109] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[5].cap_47  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net47));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[110] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[6].cap_48  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net48));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[13].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[13] ),
    .B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[111] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[13].genblk1[7].cap_49  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net49));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[112] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[0].cap_50  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net50));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[113] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[1].cap_51  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net51));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[114] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[2].cap_52  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net52));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[115] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[3].cap_53  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net53));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[116] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[4].cap_54  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net54));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[117] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[5].cap_55  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net55));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[118] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[6].cap_56  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net56));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[14].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[14] ),
    .B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[119] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[14].genblk1[7].cap_57  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net57));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[120] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[0].cap_58  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net58));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[121] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[1].cap_59  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net59));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[122] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[2].cap_60  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net60));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[123] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[3].cap_61  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net61));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[124] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[4].cap_62  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net62));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[125] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[5].cap_63  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net63));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[126] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[6].cap_64  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net64));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[15].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[15] ),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[127] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[15].genblk1[7].cap_65  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net65));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[128] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[0].cap_66  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net66));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[129] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[1].cap_67  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net67));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[130] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[2].cap_68  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net68));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[131] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[3].cap_69  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net69));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[132] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[4].cap_70  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net70));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[133] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[5].cap_71  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net71));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[134] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[6].cap_72  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net72));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[16].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[16] ),
    .B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[135] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[16].genblk1[7].cap_73  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net73));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[136] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[0].cap_74  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net74));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[137] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[1].cap_75  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net75));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[138] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[2].cap_76  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net76));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[139] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[3].cap_77  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net77));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[140] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[4].cap_78  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net78));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[141] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[5].cap_79  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net79));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[142] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[6].cap_80  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net80));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[17].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[17] ),
    .B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[143] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[17].genblk1[7].cap_81  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net81));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[144] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[0].cap_82  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net82));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[145] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[1].cap_83  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net83));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[146] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[2].cap_84  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net84));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[147] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[3].cap_85  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net85));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[148] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[4].cap_86  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net86));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[149] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[5].cap_87  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net87));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[150] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[6].cap_88  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net88));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[18].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[18] ),
    .B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[151] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[18].genblk1[7].cap_89  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net89));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[152] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[0].cap_90  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net90));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[153] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[1].cap_91  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net91));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[154] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[2].cap_92  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net92));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[155] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[3].cap_93  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net93));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[156] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[4].cap_94  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net94));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[157] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[5].cap_95  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net95));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[158] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[6].cap_96  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net96));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[19].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[19] ),
    .B(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[159] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[19].genblk1[7].cap_97  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net97));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[8] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[0].cap_98  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net98));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[9] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[1].cap_99  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net99));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[10] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[2].cap_100  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net100));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[11] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[3].cap_101  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net101));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[12] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[4].cap_102  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net102));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[13] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[5].cap_103  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net103));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[14] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[6].cap_104  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net104));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[1].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[1] ),
    .B(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[15] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[1].genblk1[7].cap_105  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net105));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[160] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[0].cap_106  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net106));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[161] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[1].cap_107  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net107));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[162] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[2].cap_108  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net108));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[163] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[3].cap_109  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net109));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[164] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[4].cap_110  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net110));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[165] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[5].cap_111  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net111));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[166] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[6].cap_112  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net112));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[20].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[20] ),
    .B(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[167] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[20].genblk1[7].cap_113  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net113));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[168] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[0].cap_114  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net114));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[169] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[1].cap_115  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net115));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[170] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[2].cap_116  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net116));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[171] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[3].cap_117  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net117));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[172] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[4].cap_118  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net118));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[173] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[5].cap_119  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net119));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[174] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[6].cap_120  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net120));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[21].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[21] ),
    .B(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[175] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[21].genblk1[7].cap_121  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net121));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[176] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[0].cap_122  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net122));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[177] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[1].cap_123  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net123));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[178] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[2].cap_124  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net124));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[179] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[3].cap_125  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net125));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[180] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[4].cap_126  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net126));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[181] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[5].cap_127  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net127));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[182] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[6].cap_128  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net128));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[22].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[22] ),
    .B(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[183] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[22].genblk1[7].cap_129  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net129));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[184] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[0].cap_130  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net130));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[185] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[1].cap_131  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net131));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[186] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[2].cap_132  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net132));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[187] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[3].cap_133  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net133));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[188] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[4].cap_134  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net134));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[189] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[5].cap_135  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net135));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[190] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[6].cap_136  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net136));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[23].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[23] ),
    .B(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[191] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[23].genblk1[7].cap_137  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net137));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[192] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[0].cap_138  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net138));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[193] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[1].cap_139  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net139));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[194] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[2].cap_140  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net140));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[195] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[3].cap_141  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net141));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[196] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[4].cap_142  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net142));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[197] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[5].cap_143  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net143));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[198] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[6].cap_144  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net144));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[24].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[24] ),
    .B(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[199] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[24].genblk1[7].cap_145  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net145));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[200] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[0].cap_146  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net146));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[201] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[1].cap_147  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net147));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[202] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[2].cap_148  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net148));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[203] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[3].cap_149  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net149));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[204] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[4].cap_150  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net150));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[205] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[5].cap_151  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net151));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[206] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[6].cap_152  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net152));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[25].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[25] ),
    .B(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[207] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[25].genblk1[7].cap_153  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net153));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[208] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[0].cap_154  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net154));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[209] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[1].cap_155  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net155));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[210] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[2].cap_156  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net156));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[211] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[3].cap_157  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net157));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[212] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[4].cap_158  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net158));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[213] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[5].cap_159  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net159));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net160),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[214] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[6].cap_160  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net160));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[26].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[26] ),
    .B(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[215] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[26].genblk1[7].cap_161  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net161));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[216] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[0].cap_162  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net162));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[217] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[1].cap_163  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net163));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net164),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[218] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[2].cap_164  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net164));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[219] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[3].cap_165  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net165));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[220] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[4].cap_166  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net166));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[221] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[5].cap_167  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net167));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[222] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[6].cap_168  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net168));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[27].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[27] ),
    .B(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[223] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[27].genblk1[7].cap_169  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net169));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[224] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[0].cap_170  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net170));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[225] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[1].cap_171  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net171));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[226] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[2].cap_172  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net172));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[227] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[3].cap_173  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net173));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[228] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[4].cap_174  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net174));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[229] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[5].cap_175  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net175));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[230] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[6].cap_176  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net176));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[28].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[28] ),
    .B(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[231] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[28].genblk1[7].cap_177  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net177));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[232] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[0].cap_178  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net178));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[233] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[1].cap_179  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net179));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[234] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[2].cap_180  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net180));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[235] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[3].cap_181  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net181));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[236] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[4].cap_182  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net182));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[237] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[5].cap_183  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net183));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[238] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[6].cap_184  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net184));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[29].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[29] ),
    .B(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[239] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[29].genblk1[7].cap_185  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net185));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[16] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[0].cap_186  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net186));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[17] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[1].cap_187  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net187));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[18] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[2].cap_188  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net188));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[19] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[3].cap_189  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net189));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[20] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[4].cap_190  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net190));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[21] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[5].cap_191  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net191));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[22] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[6].cap_192  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net192));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[2].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[2] ),
    .B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[23] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[2].genblk1[7].cap_193  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net193));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[240] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[0].cap_194  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net194));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[241] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[1].cap_195  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net195));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[242] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[2].cap_196  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net196));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[243] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[3].cap_197  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net197));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[244] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[4].cap_198  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net198));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[245] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[5].cap_199  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net199));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[246] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[6].cap_200  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net200));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[30].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[30] ),
    .B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[247] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[30].genblk1[7].cap_201  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net201));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[248] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[0].cap_202  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net202));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[249] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[1].cap_203  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net203));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[250] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[2].cap_204  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net204));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[251] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[3].cap_205  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net205));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[252] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[4].cap_206  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net206));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[253] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[5].cap_207  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net207));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[254] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[6].cap_208  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net208));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[31].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[31] ),
    .B(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[255] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[31].genblk1[7].cap_209  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net209));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[256] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[0].cap_210  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net210));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[257] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[1].cap_211  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net211));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[258] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[2].cap_212  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net212));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net213),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[259] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[3].cap_213  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net213));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[260] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[4].cap_214  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net214));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[261] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[5].cap_215  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net215));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[262] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[6].cap_216  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net216));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[32].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[32] ),
    .B(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[263] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[32].genblk1[7].cap_217  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net217));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[264] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[0].cap_218  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net218));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[265] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[1].cap_219  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net219));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[266] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[2].cap_220  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net220));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[267] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[3].cap_221  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net221));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[268] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[4].cap_222  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net222));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[269] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[5].cap_223  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net223));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[270] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[6].cap_224  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net224));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[33].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[33] ),
    .B(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[271] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[33].genblk1[7].cap_225  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net225));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[272] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[0].cap_226  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net226));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[273] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[1].cap_227  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net227));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[274] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[2].cap_228  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net228));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[275] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[3].cap_229  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net229));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[276] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[4].cap_230  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net230));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net231),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[277] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[5].cap_231  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net231));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[278] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[6].cap_232  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net232));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[34].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[34] ),
    .B(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[279] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[34].genblk1[7].cap_233  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net233));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[24] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[0].cap_234  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net234));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net235),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[25] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[1].cap_235  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net235));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[26] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[2].cap_236  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net236));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[27] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[3].cap_237  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net237));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[28] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[4].cap_238  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net238));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[29] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[5].cap_239  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net239));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[30] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[6].cap_240  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net240));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[3].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[3] ),
    .B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[31] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[3].genblk1[7].cap_241  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net241));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[32] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[0].cap_242  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net242));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[33] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[1].cap_243  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net243));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[34] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[2].cap_244  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net244));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net245),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[35] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[3].cap_245  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net245));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net246),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[36] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[4].cap_246  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net246));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[37] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[5].cap_247  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net247));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[38] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[6].cap_248  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net248));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[4].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[4] ),
    .B(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[39] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[4].genblk1[7].cap_249  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net249));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[40] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[0].cap_250  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net250));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[41] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[1].cap_251  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net251));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[42] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[2].cap_252  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net252));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[43] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[3].cap_253  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net253));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[44] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[4].cap_254  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net254));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net255),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[45] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[5].cap_255  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net255));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[46] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[6].cap_256  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net256));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[5].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[5] ),
    .B(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[47] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[5].genblk1[7].cap_257  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net257));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[48] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[0].cap_258  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net258));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[49] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[1].cap_259  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net259));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net260),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[50] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[2].cap_260  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net260));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[51] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[3].cap_261  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net261));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[52] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[4].cap_262  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net262));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[53] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[5].cap_263  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net263));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[54] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[6].cap_264  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net264));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[6].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[6] ),
    .B(net265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[55] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[6].genblk1[7].cap_265  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net265));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net266),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[56] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[0].cap_266  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net266));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net267),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[57] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[1].cap_267  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net267));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net268),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[58] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[2].cap_268  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net268));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[59] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[3].cap_269  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net269));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[60] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[4].cap_270  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net270));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net271),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[61] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[5].cap_271  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net271));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[62] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[6].cap_272  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net272));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[7].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[7] ),
    .B(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[63] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[7].genblk1[7].cap_273  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net273));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[64] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[0].cap_274  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net274));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[65] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[1].cap_275  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net275));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[66] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[2].cap_276  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net276));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[67] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[3].cap_277  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net277));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[68] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[4].cap_278  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net278));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[69] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[5].cap_279  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net279));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[70] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[6].cap_280  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net280));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[8].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[8] ),
    .B(net281),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[71] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[8].genblk1[7].cap_281  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net281));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[0].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net282),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[72] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[0].cap_282  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net282));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[1].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[73] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[1].cap_283  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net283));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[2].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net284),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[74] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[2].cap_284  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net284));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[3].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net285),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[75] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[3].cap_285  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net285));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[4].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net286),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[76] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[4].cap_286  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net286));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[5].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[77] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[5].cap_287  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net287));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[6].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net288),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[78] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[6].cap_288  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net288));
 sky130_fd_sc_hd__nand2_1 \ros_nand4_cap.genblk2[9].genblk1[7].cap  (.A(\ros_nand4_cap.nets_notouch_[9] ),
    .B(net289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\ros_nand4_cap.open_nets_notouch_[79] ));
 sky130_fd_sc_hd__conb_1 \ros_nand4_cap.genblk2[9].genblk1[7].cap_289  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net289));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net290));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net291));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net292));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net293));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net294));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net295));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net296));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net297));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net298));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net299));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net300));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net301));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net302));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net303));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net304));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net305));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net306));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net307));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net308));
 sky130_fd_sc_hd__conb_1 tt_um_gfg_development_tros_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net309));
 assign uio_oe[0] = net290;
 assign uio_oe[1] = net291;
 assign uio_oe[2] = net292;
 assign uio_oe[3] = net293;
 assign uio_oe[4] = net294;
 assign uio_oe[5] = net295;
 assign uio_oe[6] = net296;
 assign uio_oe[7] = net297;
 assign uio_out[0] = net298;
 assign uio_out[1] = net299;
 assign uio_out[2] = net300;
 assign uio_out[3] = net301;
 assign uio_out[4] = net302;
 assign uio_out[5] = net303;
 assign uio_out[6] = net304;
 assign uio_out[7] = net305;
 assign uo_out[0] = net306;
 assign uo_out[1] = net307;
 assign uo_out[2] = net308;
 assign uo_out[3] = net309;
endmodule
